module vsdbabysoc (ENb_CP,
    ENb_VCO,
    OUT,
    REF,
    VCO_IN,
    VREFH,
    reset);
 input ENb_CP;
 input ENb_VCO;
 output OUT;
 input REF;
 input VCO_IN;
 input VREFH;
 input reset;

 wire CLK;
 wire net10;
 wire \RV_TO_DAC[0] ;
 wire \RV_TO_DAC[1] ;
 wire \RV_TO_DAC[2] ;
 wire \RV_TO_DAC[3] ;
 wire \RV_TO_DAC[4] ;
 wire \RV_TO_DAC[5] ;
 wire \RV_TO_DAC[6] ;
 wire \RV_TO_DAC[7] ;
 wire \RV_TO_DAC[8] ;
 wire \RV_TO_DAC[9] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01122_;
 wire _01127_;
 wire _01130_;
 wire _01133_;
 wire _01136_;
 wire _01137_;
 wire _01142_;
 wire _01146_;
 wire _01151_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01157_;
 wire _01159_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01170_;
 wire _01176_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01191_;
 wire _01195_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01202_;
 wire _01203_;
 wire _01206_;
 wire _01207_;
 wire _01209_;
 wire _01215_;
 wire _01216_;
 wire _01219_;
 wire _01220_;
 wire _01223_;
 wire _01224_;
 wire _01227_;
 wire _01228_;
 wire _01231_;
 wire _01232_;
 wire _01235_;
 wire _01236_;
 wire _01239_;
 wire _01240_;
 wire _01243_;
 wire _01244_;
 wire _01247_;
 wire _01248_;
 wire _01252_;
 wire _01254_;
 wire _01258_;
 wire _01259_;
 wire _01262_;
 wire _01263_;
 wire _01266_;
 wire _01267_;
 wire _01270_;
 wire _01271_;
 wire _01274_;
 wire _01275_;
 wire _01278_;
 wire _01279_;
 wire _01282_;
 wire _01283_;
 wire _01286_;
 wire _01287_;
 wire _01290_;
 wire _01291_;
 wire _01295_;
 wire _01297_;
 wire _01301_;
 wire _01302_;
 wire _01305_;
 wire _01306_;
 wire _01309_;
 wire _01310_;
 wire _01313_;
 wire _01314_;
 wire _01317_;
 wire _01318_;
 wire _01321_;
 wire _01322_;
 wire _01325_;
 wire _01326_;
 wire _01329_;
 wire _01330_;
 wire _01333_;
 wire _01334_;
 wire _01337_;
 wire _01338_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01346_;
 wire _01348_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01370_;
 wire _01372_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01396_;
 wire _01398_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01429_;
 wire _01430_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01448_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01473_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01503_;
 wire _01504_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01526_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01549_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01580_;
 wire _01582_;
 wire _01583_;
 wire _01585_;
 wire _01586_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01604_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01627_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01663_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01678_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01704_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01737_;
 wire _01738_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire clknet_4_15_0_CLK;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire clknet_4_14_0_CLK;
 wire _01756_;
 wire clknet_4_13_0_CLK;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire clknet_4_12_0_CLK;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire clknet_4_11_0_CLK;
 wire _01781_;
 wire clknet_4_10_0_CLK;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire clknet_4_9_0_CLK;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire clknet_4_8_0_CLK;
 wire _01813_;
 wire clknet_4_7_0_CLK;
 wire _01815_;
 wire _01816_;
 wire clknet_4_6_0_CLK;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire clknet_4_5_0_CLK;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire clknet_4_4_0_CLK;
 wire _01839_;
 wire clknet_4_3_0_CLK;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire clknet_4_2_0_CLK;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire clknet_4_1_0_CLK;
 wire _01862_;
 wire clknet_4_0_0_CLK;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire clknet_0_CLK;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire clknet_leaf_112_CLK;
 wire _01890_;
 wire _01891_;
 wire clknet_leaf_111_CLK;
 wire _01893_;
 wire clknet_leaf_110_CLK;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire clknet_leaf_109_CLK;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire clknet_leaf_108_CLK;
 wire _01914_;
 wire clknet_leaf_107_CLK;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire clknet_leaf_106_CLK;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire clknet_leaf_105_CLK;
 wire _01939_;
 wire clknet_leaf_104_CLK;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire clknet_leaf_103_CLK;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire clknet_leaf_102_CLK;
 wire _01967_;
 wire clknet_leaf_101_CLK;
 wire _01969_;
 wire _01970_;
 wire clknet_leaf_100_CLK;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire clknet_leaf_99_CLK;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire clknet_leaf_98_CLK;
 wire _01991_;
 wire clknet_leaf_97_CLK;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire clknet_leaf_96_CLK;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire clknet_leaf_95_CLK;
 wire clknet_leaf_94_CLK;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire clknet_leaf_93_CLK;
 wire _02018_;
 wire clknet_leaf_92_CLK;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire clknet_leaf_91_CLK;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire clknet_leaf_90_CLK;
 wire _02046_;
 wire clknet_leaf_89_CLK;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire clknet_leaf_88_CLK;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire clknet_leaf_87_CLK;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire clknet_leaf_86_CLK;
 wire _02071_;
 wire clknet_leaf_85_CLK;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire clknet_leaf_84_CLK;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire clknet_leaf_83_CLK;
 wire _02094_;
 wire clknet_leaf_82_CLK;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire clknet_leaf_81_CLK;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire clknet_leaf_80_CLK;
 wire _02125_;
 wire _02126_;
 wire clknet_leaf_79_CLK;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire clknet_leaf_78_CLK;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire clknet_leaf_77_CLK;
 wire _02147_;
 wire clknet_leaf_76_CLK;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire clknet_leaf_75_CLK;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire clknet_leaf_74_CLK;
 wire _02170_;
 wire clknet_leaf_73_CLK;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire clknet_leaf_72_CLK;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire clknet_leaf_71_CLK;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire clknet_leaf_70_CLK;
 wire _02204_;
 wire clknet_leaf_69_CLK;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire clknet_leaf_68_CLK;
 wire _02221_;
 wire clknet_leaf_67_CLK;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire clknet_leaf_66_CLK;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire clknet_leaf_65_CLK;
 wire _02246_;
 wire clknet_leaf_64_CLK;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire clknet_leaf_63_CLK;
 wire clknet_leaf_62_CLK;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire clknet_leaf_61_CLK;
 wire _02277_;
 wire clknet_leaf_60_CLK;
 wire _02279_;
 wire _02280_;
 wire clknet_leaf_59_CLK;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire clknet_leaf_58_CLK;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire clknet_leaf_57_CLK;
 wire _02299_;
 wire clknet_leaf_56_CLK;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire clknet_leaf_55_CLK;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire clknet_leaf_54_CLK;
 wire _02324_;
 wire clknet_leaf_53_CLK;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire clknet_leaf_52_CLK;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire clknet_leaf_51_CLK;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire clknet_leaf_50_CLK;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire clknet_leaf_49_CLK;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire clknet_leaf_48_CLK;
 wire _02377_;
 wire clknet_leaf_47_CLK;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire clknet_leaf_46_CLK;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire clknet_leaf_45_CLK;
 wire _02400_;
 wire clknet_leaf_44_CLK;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire clknet_leaf_43_CLK;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire clknet_leaf_42_CLK;
 wire _02430_;
 wire clknet_leaf_41_CLK;
 wire _02432_;
 wire _02433_;
 wire clknet_leaf_40_CLK;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire clknet_leaf_39_CLK;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire clknet_leaf_38_CLK;
 wire _02454_;
 wire clknet_leaf_37_CLK;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire clknet_leaf_36_CLK;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire clknet_leaf_35_CLK;
 wire _02477_;
 wire clknet_leaf_34_CLK;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire clknet_leaf_33_CLK;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire clknet_leaf_32_CLK;
 wire clknet_leaf_31_CLK;
 wire clknet_leaf_30_CLK;
 wire clknet_leaf_29_CLK;
 wire clknet_leaf_28_CLK;
 wire clknet_leaf_27_CLK;
 wire clknet_leaf_26_CLK;
 wire _02512_;
 wire clknet_leaf_25_CLK;
 wire clknet_leaf_24_CLK;
 wire clknet_leaf_23_CLK;
 wire clknet_leaf_22_CLK;
 wire _02517_;
 wire clknet_leaf_21_CLK;
 wire clknet_leaf_20_CLK;
 wire clknet_leaf_19_CLK;
 wire _02521_;
 wire clknet_leaf_18_CLK;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire clknet_leaf_17_CLK;
 wire _02527_;
 wire _02528_;
 wire clknet_leaf_16_CLK;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire clknet_leaf_15_CLK;
 wire _02539_;
 wire _02540_;
 wire clknet_leaf_14_CLK;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire clknet_leaf_13_CLK;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire clknet_leaf_12_CLK;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire clknet_leaf_11_CLK;
 wire clknet_leaf_10_CLK;
 wire _02566_;
 wire clknet_leaf_9_CLK;
 wire clknet_leaf_8_CLK;
 wire clknet_leaf_7_CLK;
 wire _02570_;
 wire clknet_leaf_6_CLK;
 wire _02572_;
 wire _02573_;
 wire clknet_leaf_5_CLK;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire clknet_leaf_4_CLK;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire net605;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire net604;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire net603;
 wire _02644_;
 wire net602;
 wire net601;
 wire net596;
 wire net594;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire net592;
 wire _02721_;
 wire net590;
 wire net588;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire net587;
 wire _02728_;
 wire _02729_;
 wire net586;
 wire net585;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire net584;
 wire _02741_;
 wire net583;
 wire _02743_;
 wire net582;
 wire _02745_;
 wire net581;
 wire _02747_;
 wire _02748_;
 wire net580;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire net579;
 wire net578;
 wire _02763_;
 wire _02764_;
 wire net577;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire net576;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire net575;
 wire net574;
 wire _02814_;
 wire net573;
 wire net572;
 wire net571;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire net570;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire net569;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire net568;
 wire net567;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire net566;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire net565;
 wire _02956_;
 wire _02957_;
 wire net564;
 wire net559;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire net558;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire net552;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire net551;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire net550;
 wire net548;
 wire _03006_;
 wire net545;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire net542;
 wire net541;
 wire _03046_;
 wire net540;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire net539;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire net536;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire net532;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire net530;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire net528;
 wire _03311_;
 wire net524;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire net520;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire net516;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire net512;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire net510;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire net508;
 wire net506;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire net504;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire net502;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire net500;
 wire _03539_;
 wire net498;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire net496;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire net494;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire net492;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire net489;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire net487;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire net480;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire net478;
 wire net472;
 wire net470;
 wire _03755_;
 wire net469;
 wire _03757_;
 wire _03758_;
 wire net468;
 wire _03760_;
 wire _03761_;
 wire net466;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire net483;
 wire _03768_;
 wire net485;
 wire net482;
 wire _03771_;
 wire net481;
 wire _03773_;
 wire _03774_;
 wire net479;
 wire net477;
 wire _03777_;
 wire net476;
 wire _03779_;
 wire net475;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire net473;
 wire _03786_;
 wire net474;
 wire _03788_;
 wire _03789_;
 wire net471;
 wire _03791_;
 wire net467;
 wire _03793_;
 wire net463;
 wire _03795_;
 wire _03796_;
 wire net443;
 wire _03798_;
 wire _03799_;
 wire net430;
 wire net429;
 wire _03802_;
 wire _03803_;
 wire net428;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire net425;
 wire net424;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire net423;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire net420;
 wire _03820_;
 wire net419;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire net417;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire net412;
 wire net410;
 wire _03839_;
 wire net408;
 wire net406;
 wire _03842_;
 wire _03843_;
 wire net403;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire net395;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire net393;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire net392;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire net391;
 wire net394;
 wire net390;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire net378;
 wire _03903_;
 wire net376;
 wire _03905_;
 wire net375;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire net374;
 wire net379;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire net372;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire net370;
 wire net371;
 wire net369;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire net367;
 wire net365;
 wire net364;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire net363;
 wire _03965_;
 wire net361;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire net360;
 wire net357;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire net356;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire net355;
 wire net354;
 wire net353;
 wire net348;
 wire _04018_;
 wire net347;
 wire _04020_;
 wire _04021_;
 wire net346;
 wire _04023_;
 wire net345;
 wire net611;
 wire _04026_;
 wire _04027_;
 wire net610;
 wire _04029_;
 wire net612;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire net608;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire net609;
 wire net613;
 wire clknet_leaf_1_CLK;
 wire _04075_;
 wire net599;
 wire net600;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire net598;
 wire _04082_;
 wire _04083_;
 wire net595;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire net593;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire net591;
 wire _04126_;
 wire _04127_;
 wire net589;
 wire _04129_;
 wire net563;
 wire net597;
 wire _04132_;
 wire net561;
 wire _04134_;
 wire net562;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire net560;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire net555;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire net554;
 wire net556;
 wire net538;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire net537;
 wire _04190_;
 wire net535;
 wire _04192_;
 wire _04193_;
 wire net543;
 wire _04195_;
 wire _04196_;
 wire net534;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire net544;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire net533;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire net531;
 wire _04239_;
 wire _04240_;
 wire net546;
 wire _04242_;
 wire net529;
 wire net547;
 wire _04245_;
 wire _04246_;
 wire net557;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire net553;
 wire clknet_leaf_2_CLK;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire net527;
 wire net549;
 wire net607;
 wire _04294_;
 wire _04295_;
 wire clknet_leaf_3_CLK;
 wire _04297_;
 wire _04298_;
 wire net526;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire net525;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire net606;
 wire _04393_;
 wire _04394_;
 wire net523;
 wire _04396_;
 wire net614;
 wire _04398_;
 wire _04399_;
 wire net615;
 wire net522;
 wire clknet_leaf_0_CLK;
 wire net521;
 wire net519;
 wire net620;
 wire _04406_;
 wire net619;
 wire net518;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire net617;
 wire _04415_;
 wire _04416_;
 wire net618;
 wire net517;
 wire _04419_;
 wire net381;
 wire net382;
 wire _04422_;
 wire net349;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire net515;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire net616;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire net404;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire net387;
 wire _04445_;
 wire _04446_;
 wire net513;
 wire net409;
 wire net514;
 wire net350;
 wire _04451_;
 wire _04452_;
 wire net344;
 wire net511;
 wire _04455_;
 wire net368;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire net509;
 wire _04462_;
 wire net351;
 wire _04464_;
 wire net385;
 wire _04466_;
 wire _04467_;
 wire net383;
 wire _04469_;
 wire net507;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire net380;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire net384;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire net386;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire net388;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire net389;
 wire net505;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire net503;
 wire net396;
 wire _04748_;
 wire net397;
 wire net501;
 wire _04751_;
 wire _04752_;
 wire net398;
 wire net499;
 wire _04755_;
 wire net399;
 wire net400;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire net401;
 wire _04762_;
 wire _04763_;
 wire net497;
 wire net495;
 wire net493;
 wire net402;
 wire net405;
 wire net491;
 wire net407;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire net433;
 wire _04776_;
 wire net434;
 wire net490;
 wire _04779_;
 wire net460;
 wire net488;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire net459;
 wire _04786_;
 wire net461;
 wire _04788_;
 wire net486;
 wire net464;
 wire _04791_;
 wire net465;
 wire _04793_;
 wire _04794_;
 wire net484;
 wire net462;
 wire _04797_;
 wire net458;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire net457;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire net456;
 wire _04808_;
 wire net455;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire net454;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire net453;
 wire net452;
 wire net451;
 wire _05030_;
 wire net450;
 wire net449;
 wire _05033_;
 wire net448;
 wire net447;
 wire _05036_;
 wire net446;
 wire net445;
 wire _05039_;
 wire _05040_;
 wire net444;
 wire net440;
 wire _05043_;
 wire net439;
 wire net442;
 wire _05046_;
 wire net438;
 wire net437;
 wire _05049_;
 wire net435;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire net441;
 wire net436;
 wire _05056_;
 wire net432;
 wire _05058_;
 wire net427;
 wire _05060_;
 wire _05061_;
 wire net431;
 wire net426;
 wire _05064_;
 wire _05065_;
 wire net422;
 wire net421;
 wire _05068_;
 wire net418;
 wire _05070_;
 wire _05071_;
 wire net416;
 wire _05073_;
 wire net414;
 wire _05075_;
 wire net413;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire net415;
 wire net411;
 wire _05083_;
 wire net377;
 wire _05085_;
 wire net373;
 wire _05087_;
 wire _05088_;
 wire net366;
 wire _05090_;
 wire net359;
 wire _05092_;
 wire _05093_;
 wire net358;
 wire _05095_;
 wire _05096_;
 wire net362;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire net352;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire net9;
 wire _05137_;
 wire _05138_;
 wire net8;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire net7;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire net6;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire net5;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire net4;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire \core.CPU_Dmem_value_a5[0][0] ;
 wire \core.CPU_Dmem_value_a5[0][10] ;
 wire \core.CPU_Dmem_value_a5[0][11] ;
 wire \core.CPU_Dmem_value_a5[0][12] ;
 wire \core.CPU_Dmem_value_a5[0][13] ;
 wire \core.CPU_Dmem_value_a5[0][14] ;
 wire \core.CPU_Dmem_value_a5[0][15] ;
 wire \core.CPU_Dmem_value_a5[0][16] ;
 wire \core.CPU_Dmem_value_a5[0][17] ;
 wire \core.CPU_Dmem_value_a5[0][18] ;
 wire \core.CPU_Dmem_value_a5[0][19] ;
 wire \core.CPU_Dmem_value_a5[0][1] ;
 wire \core.CPU_Dmem_value_a5[0][20] ;
 wire \core.CPU_Dmem_value_a5[0][21] ;
 wire \core.CPU_Dmem_value_a5[0][22] ;
 wire \core.CPU_Dmem_value_a5[0][23] ;
 wire \core.CPU_Dmem_value_a5[0][24] ;
 wire \core.CPU_Dmem_value_a5[0][25] ;
 wire \core.CPU_Dmem_value_a5[0][26] ;
 wire \core.CPU_Dmem_value_a5[0][27] ;
 wire \core.CPU_Dmem_value_a5[0][28] ;
 wire \core.CPU_Dmem_value_a5[0][29] ;
 wire \core.CPU_Dmem_value_a5[0][2] ;
 wire \core.CPU_Dmem_value_a5[0][30] ;
 wire \core.CPU_Dmem_value_a5[0][31] ;
 wire \core.CPU_Dmem_value_a5[0][3] ;
 wire \core.CPU_Dmem_value_a5[0][4] ;
 wire \core.CPU_Dmem_value_a5[0][5] ;
 wire \core.CPU_Dmem_value_a5[0][6] ;
 wire \core.CPU_Dmem_value_a5[0][7] ;
 wire \core.CPU_Dmem_value_a5[0][8] ;
 wire \core.CPU_Dmem_value_a5[0][9] ;
 wire \core.CPU_Dmem_value_a5[10][0] ;
 wire \core.CPU_Dmem_value_a5[10][10] ;
 wire \core.CPU_Dmem_value_a5[10][11] ;
 wire \core.CPU_Dmem_value_a5[10][12] ;
 wire \core.CPU_Dmem_value_a5[10][13] ;
 wire \core.CPU_Dmem_value_a5[10][14] ;
 wire \core.CPU_Dmem_value_a5[10][15] ;
 wire \core.CPU_Dmem_value_a5[10][16] ;
 wire \core.CPU_Dmem_value_a5[10][17] ;
 wire \core.CPU_Dmem_value_a5[10][18] ;
 wire \core.CPU_Dmem_value_a5[10][19] ;
 wire \core.CPU_Dmem_value_a5[10][1] ;
 wire \core.CPU_Dmem_value_a5[10][20] ;
 wire \core.CPU_Dmem_value_a5[10][21] ;
 wire \core.CPU_Dmem_value_a5[10][22] ;
 wire \core.CPU_Dmem_value_a5[10][23] ;
 wire \core.CPU_Dmem_value_a5[10][24] ;
 wire \core.CPU_Dmem_value_a5[10][25] ;
 wire \core.CPU_Dmem_value_a5[10][26] ;
 wire \core.CPU_Dmem_value_a5[10][27] ;
 wire \core.CPU_Dmem_value_a5[10][28] ;
 wire \core.CPU_Dmem_value_a5[10][29] ;
 wire \core.CPU_Dmem_value_a5[10][2] ;
 wire \core.CPU_Dmem_value_a5[10][30] ;
 wire \core.CPU_Dmem_value_a5[10][31] ;
 wire \core.CPU_Dmem_value_a5[10][3] ;
 wire \core.CPU_Dmem_value_a5[10][4] ;
 wire \core.CPU_Dmem_value_a5[10][5] ;
 wire \core.CPU_Dmem_value_a5[10][6] ;
 wire \core.CPU_Dmem_value_a5[10][7] ;
 wire \core.CPU_Dmem_value_a5[10][8] ;
 wire \core.CPU_Dmem_value_a5[10][9] ;
 wire \core.CPU_Dmem_value_a5[11][0] ;
 wire \core.CPU_Dmem_value_a5[11][10] ;
 wire \core.CPU_Dmem_value_a5[11][11] ;
 wire \core.CPU_Dmem_value_a5[11][12] ;
 wire \core.CPU_Dmem_value_a5[11][13] ;
 wire \core.CPU_Dmem_value_a5[11][14] ;
 wire \core.CPU_Dmem_value_a5[11][15] ;
 wire \core.CPU_Dmem_value_a5[11][16] ;
 wire \core.CPU_Dmem_value_a5[11][17] ;
 wire \core.CPU_Dmem_value_a5[11][18] ;
 wire \core.CPU_Dmem_value_a5[11][19] ;
 wire \core.CPU_Dmem_value_a5[11][1] ;
 wire \core.CPU_Dmem_value_a5[11][20] ;
 wire \core.CPU_Dmem_value_a5[11][21] ;
 wire \core.CPU_Dmem_value_a5[11][22] ;
 wire \core.CPU_Dmem_value_a5[11][23] ;
 wire \core.CPU_Dmem_value_a5[11][24] ;
 wire \core.CPU_Dmem_value_a5[11][25] ;
 wire \core.CPU_Dmem_value_a5[11][26] ;
 wire \core.CPU_Dmem_value_a5[11][27] ;
 wire \core.CPU_Dmem_value_a5[11][28] ;
 wire \core.CPU_Dmem_value_a5[11][29] ;
 wire \core.CPU_Dmem_value_a5[11][2] ;
 wire \core.CPU_Dmem_value_a5[11][30] ;
 wire \core.CPU_Dmem_value_a5[11][31] ;
 wire \core.CPU_Dmem_value_a5[11][3] ;
 wire \core.CPU_Dmem_value_a5[11][4] ;
 wire \core.CPU_Dmem_value_a5[11][5] ;
 wire \core.CPU_Dmem_value_a5[11][6] ;
 wire \core.CPU_Dmem_value_a5[11][7] ;
 wire \core.CPU_Dmem_value_a5[11][8] ;
 wire \core.CPU_Dmem_value_a5[11][9] ;
 wire \core.CPU_Dmem_value_a5[12][0] ;
 wire \core.CPU_Dmem_value_a5[12][10] ;
 wire \core.CPU_Dmem_value_a5[12][11] ;
 wire \core.CPU_Dmem_value_a5[12][12] ;
 wire \core.CPU_Dmem_value_a5[12][13] ;
 wire \core.CPU_Dmem_value_a5[12][14] ;
 wire \core.CPU_Dmem_value_a5[12][15] ;
 wire \core.CPU_Dmem_value_a5[12][16] ;
 wire \core.CPU_Dmem_value_a5[12][17] ;
 wire \core.CPU_Dmem_value_a5[12][18] ;
 wire \core.CPU_Dmem_value_a5[12][19] ;
 wire \core.CPU_Dmem_value_a5[12][1] ;
 wire \core.CPU_Dmem_value_a5[12][20] ;
 wire \core.CPU_Dmem_value_a5[12][21] ;
 wire \core.CPU_Dmem_value_a5[12][22] ;
 wire \core.CPU_Dmem_value_a5[12][23] ;
 wire \core.CPU_Dmem_value_a5[12][24] ;
 wire \core.CPU_Dmem_value_a5[12][25] ;
 wire \core.CPU_Dmem_value_a5[12][26] ;
 wire \core.CPU_Dmem_value_a5[12][27] ;
 wire \core.CPU_Dmem_value_a5[12][28] ;
 wire \core.CPU_Dmem_value_a5[12][29] ;
 wire \core.CPU_Dmem_value_a5[12][2] ;
 wire \core.CPU_Dmem_value_a5[12][30] ;
 wire \core.CPU_Dmem_value_a5[12][31] ;
 wire \core.CPU_Dmem_value_a5[12][3] ;
 wire \core.CPU_Dmem_value_a5[12][4] ;
 wire \core.CPU_Dmem_value_a5[12][5] ;
 wire \core.CPU_Dmem_value_a5[12][6] ;
 wire \core.CPU_Dmem_value_a5[12][7] ;
 wire \core.CPU_Dmem_value_a5[12][8] ;
 wire \core.CPU_Dmem_value_a5[12][9] ;
 wire \core.CPU_Dmem_value_a5[13][0] ;
 wire \core.CPU_Dmem_value_a5[13][10] ;
 wire \core.CPU_Dmem_value_a5[13][11] ;
 wire \core.CPU_Dmem_value_a5[13][12] ;
 wire \core.CPU_Dmem_value_a5[13][13] ;
 wire \core.CPU_Dmem_value_a5[13][14] ;
 wire \core.CPU_Dmem_value_a5[13][15] ;
 wire \core.CPU_Dmem_value_a5[13][16] ;
 wire \core.CPU_Dmem_value_a5[13][17] ;
 wire \core.CPU_Dmem_value_a5[13][18] ;
 wire \core.CPU_Dmem_value_a5[13][19] ;
 wire \core.CPU_Dmem_value_a5[13][1] ;
 wire \core.CPU_Dmem_value_a5[13][20] ;
 wire \core.CPU_Dmem_value_a5[13][21] ;
 wire \core.CPU_Dmem_value_a5[13][22] ;
 wire \core.CPU_Dmem_value_a5[13][23] ;
 wire \core.CPU_Dmem_value_a5[13][24] ;
 wire \core.CPU_Dmem_value_a5[13][25] ;
 wire \core.CPU_Dmem_value_a5[13][26] ;
 wire \core.CPU_Dmem_value_a5[13][27] ;
 wire \core.CPU_Dmem_value_a5[13][28] ;
 wire \core.CPU_Dmem_value_a5[13][29] ;
 wire \core.CPU_Dmem_value_a5[13][2] ;
 wire \core.CPU_Dmem_value_a5[13][30] ;
 wire \core.CPU_Dmem_value_a5[13][31] ;
 wire \core.CPU_Dmem_value_a5[13][3] ;
 wire \core.CPU_Dmem_value_a5[13][4] ;
 wire \core.CPU_Dmem_value_a5[13][5] ;
 wire \core.CPU_Dmem_value_a5[13][6] ;
 wire \core.CPU_Dmem_value_a5[13][7] ;
 wire \core.CPU_Dmem_value_a5[13][8] ;
 wire \core.CPU_Dmem_value_a5[13][9] ;
 wire \core.CPU_Dmem_value_a5[14][0] ;
 wire \core.CPU_Dmem_value_a5[14][10] ;
 wire \core.CPU_Dmem_value_a5[14][11] ;
 wire \core.CPU_Dmem_value_a5[14][12] ;
 wire \core.CPU_Dmem_value_a5[14][13] ;
 wire \core.CPU_Dmem_value_a5[14][14] ;
 wire \core.CPU_Dmem_value_a5[14][15] ;
 wire \core.CPU_Dmem_value_a5[14][16] ;
 wire \core.CPU_Dmem_value_a5[14][17] ;
 wire \core.CPU_Dmem_value_a5[14][18] ;
 wire \core.CPU_Dmem_value_a5[14][19] ;
 wire \core.CPU_Dmem_value_a5[14][1] ;
 wire \core.CPU_Dmem_value_a5[14][20] ;
 wire \core.CPU_Dmem_value_a5[14][21] ;
 wire \core.CPU_Dmem_value_a5[14][22] ;
 wire \core.CPU_Dmem_value_a5[14][23] ;
 wire \core.CPU_Dmem_value_a5[14][24] ;
 wire \core.CPU_Dmem_value_a5[14][25] ;
 wire \core.CPU_Dmem_value_a5[14][26] ;
 wire \core.CPU_Dmem_value_a5[14][27] ;
 wire \core.CPU_Dmem_value_a5[14][28] ;
 wire \core.CPU_Dmem_value_a5[14][29] ;
 wire \core.CPU_Dmem_value_a5[14][2] ;
 wire \core.CPU_Dmem_value_a5[14][30] ;
 wire \core.CPU_Dmem_value_a5[14][31] ;
 wire \core.CPU_Dmem_value_a5[14][3] ;
 wire \core.CPU_Dmem_value_a5[14][4] ;
 wire \core.CPU_Dmem_value_a5[14][5] ;
 wire \core.CPU_Dmem_value_a5[14][6] ;
 wire \core.CPU_Dmem_value_a5[14][7] ;
 wire \core.CPU_Dmem_value_a5[14][8] ;
 wire \core.CPU_Dmem_value_a5[14][9] ;
 wire \core.CPU_Dmem_value_a5[15][0] ;
 wire \core.CPU_Dmem_value_a5[15][10] ;
 wire \core.CPU_Dmem_value_a5[15][11] ;
 wire \core.CPU_Dmem_value_a5[15][12] ;
 wire \core.CPU_Dmem_value_a5[15][13] ;
 wire \core.CPU_Dmem_value_a5[15][14] ;
 wire \core.CPU_Dmem_value_a5[15][15] ;
 wire \core.CPU_Dmem_value_a5[15][16] ;
 wire \core.CPU_Dmem_value_a5[15][17] ;
 wire \core.CPU_Dmem_value_a5[15][18] ;
 wire \core.CPU_Dmem_value_a5[15][19] ;
 wire \core.CPU_Dmem_value_a5[15][1] ;
 wire \core.CPU_Dmem_value_a5[15][20] ;
 wire \core.CPU_Dmem_value_a5[15][21] ;
 wire \core.CPU_Dmem_value_a5[15][22] ;
 wire \core.CPU_Dmem_value_a5[15][23] ;
 wire \core.CPU_Dmem_value_a5[15][24] ;
 wire \core.CPU_Dmem_value_a5[15][25] ;
 wire \core.CPU_Dmem_value_a5[15][26] ;
 wire \core.CPU_Dmem_value_a5[15][27] ;
 wire \core.CPU_Dmem_value_a5[15][28] ;
 wire \core.CPU_Dmem_value_a5[15][29] ;
 wire \core.CPU_Dmem_value_a5[15][2] ;
 wire \core.CPU_Dmem_value_a5[15][30] ;
 wire \core.CPU_Dmem_value_a5[15][31] ;
 wire \core.CPU_Dmem_value_a5[15][3] ;
 wire \core.CPU_Dmem_value_a5[15][4] ;
 wire \core.CPU_Dmem_value_a5[15][5] ;
 wire \core.CPU_Dmem_value_a5[15][6] ;
 wire \core.CPU_Dmem_value_a5[15][7] ;
 wire \core.CPU_Dmem_value_a5[15][8] ;
 wire \core.CPU_Dmem_value_a5[15][9] ;
 wire \core.CPU_Dmem_value_a5[1][0] ;
 wire \core.CPU_Dmem_value_a5[1][10] ;
 wire \core.CPU_Dmem_value_a5[1][11] ;
 wire \core.CPU_Dmem_value_a5[1][12] ;
 wire \core.CPU_Dmem_value_a5[1][13] ;
 wire \core.CPU_Dmem_value_a5[1][14] ;
 wire \core.CPU_Dmem_value_a5[1][15] ;
 wire \core.CPU_Dmem_value_a5[1][16] ;
 wire \core.CPU_Dmem_value_a5[1][17] ;
 wire \core.CPU_Dmem_value_a5[1][18] ;
 wire \core.CPU_Dmem_value_a5[1][19] ;
 wire \core.CPU_Dmem_value_a5[1][1] ;
 wire \core.CPU_Dmem_value_a5[1][20] ;
 wire \core.CPU_Dmem_value_a5[1][21] ;
 wire \core.CPU_Dmem_value_a5[1][22] ;
 wire \core.CPU_Dmem_value_a5[1][23] ;
 wire \core.CPU_Dmem_value_a5[1][24] ;
 wire \core.CPU_Dmem_value_a5[1][25] ;
 wire \core.CPU_Dmem_value_a5[1][26] ;
 wire \core.CPU_Dmem_value_a5[1][27] ;
 wire \core.CPU_Dmem_value_a5[1][28] ;
 wire \core.CPU_Dmem_value_a5[1][29] ;
 wire \core.CPU_Dmem_value_a5[1][2] ;
 wire \core.CPU_Dmem_value_a5[1][30] ;
 wire \core.CPU_Dmem_value_a5[1][31] ;
 wire \core.CPU_Dmem_value_a5[1][3] ;
 wire \core.CPU_Dmem_value_a5[1][4] ;
 wire \core.CPU_Dmem_value_a5[1][5] ;
 wire \core.CPU_Dmem_value_a5[1][6] ;
 wire \core.CPU_Dmem_value_a5[1][7] ;
 wire \core.CPU_Dmem_value_a5[1][8] ;
 wire \core.CPU_Dmem_value_a5[1][9] ;
 wire \core.CPU_Dmem_value_a5[2][0] ;
 wire \core.CPU_Dmem_value_a5[2][10] ;
 wire \core.CPU_Dmem_value_a5[2][11] ;
 wire \core.CPU_Dmem_value_a5[2][12] ;
 wire \core.CPU_Dmem_value_a5[2][13] ;
 wire \core.CPU_Dmem_value_a5[2][14] ;
 wire \core.CPU_Dmem_value_a5[2][15] ;
 wire \core.CPU_Dmem_value_a5[2][16] ;
 wire \core.CPU_Dmem_value_a5[2][17] ;
 wire \core.CPU_Dmem_value_a5[2][18] ;
 wire \core.CPU_Dmem_value_a5[2][19] ;
 wire \core.CPU_Dmem_value_a5[2][1] ;
 wire \core.CPU_Dmem_value_a5[2][20] ;
 wire \core.CPU_Dmem_value_a5[2][21] ;
 wire \core.CPU_Dmem_value_a5[2][22] ;
 wire \core.CPU_Dmem_value_a5[2][23] ;
 wire \core.CPU_Dmem_value_a5[2][24] ;
 wire \core.CPU_Dmem_value_a5[2][25] ;
 wire \core.CPU_Dmem_value_a5[2][26] ;
 wire \core.CPU_Dmem_value_a5[2][27] ;
 wire \core.CPU_Dmem_value_a5[2][28] ;
 wire \core.CPU_Dmem_value_a5[2][29] ;
 wire \core.CPU_Dmem_value_a5[2][2] ;
 wire \core.CPU_Dmem_value_a5[2][30] ;
 wire \core.CPU_Dmem_value_a5[2][31] ;
 wire \core.CPU_Dmem_value_a5[2][3] ;
 wire \core.CPU_Dmem_value_a5[2][4] ;
 wire \core.CPU_Dmem_value_a5[2][5] ;
 wire \core.CPU_Dmem_value_a5[2][6] ;
 wire \core.CPU_Dmem_value_a5[2][7] ;
 wire \core.CPU_Dmem_value_a5[2][8] ;
 wire \core.CPU_Dmem_value_a5[2][9] ;
 wire \core.CPU_Dmem_value_a5[3][0] ;
 wire \core.CPU_Dmem_value_a5[3][10] ;
 wire \core.CPU_Dmem_value_a5[3][11] ;
 wire \core.CPU_Dmem_value_a5[3][12] ;
 wire \core.CPU_Dmem_value_a5[3][13] ;
 wire \core.CPU_Dmem_value_a5[3][14] ;
 wire \core.CPU_Dmem_value_a5[3][15] ;
 wire \core.CPU_Dmem_value_a5[3][16] ;
 wire \core.CPU_Dmem_value_a5[3][17] ;
 wire \core.CPU_Dmem_value_a5[3][18] ;
 wire \core.CPU_Dmem_value_a5[3][19] ;
 wire \core.CPU_Dmem_value_a5[3][1] ;
 wire \core.CPU_Dmem_value_a5[3][20] ;
 wire \core.CPU_Dmem_value_a5[3][21] ;
 wire \core.CPU_Dmem_value_a5[3][22] ;
 wire \core.CPU_Dmem_value_a5[3][23] ;
 wire \core.CPU_Dmem_value_a5[3][24] ;
 wire \core.CPU_Dmem_value_a5[3][25] ;
 wire \core.CPU_Dmem_value_a5[3][26] ;
 wire \core.CPU_Dmem_value_a5[3][27] ;
 wire \core.CPU_Dmem_value_a5[3][28] ;
 wire \core.CPU_Dmem_value_a5[3][29] ;
 wire \core.CPU_Dmem_value_a5[3][2] ;
 wire \core.CPU_Dmem_value_a5[3][30] ;
 wire \core.CPU_Dmem_value_a5[3][31] ;
 wire \core.CPU_Dmem_value_a5[3][3] ;
 wire \core.CPU_Dmem_value_a5[3][4] ;
 wire \core.CPU_Dmem_value_a5[3][5] ;
 wire \core.CPU_Dmem_value_a5[3][6] ;
 wire \core.CPU_Dmem_value_a5[3][7] ;
 wire \core.CPU_Dmem_value_a5[3][8] ;
 wire \core.CPU_Dmem_value_a5[3][9] ;
 wire \core.CPU_Dmem_value_a5[4][0] ;
 wire \core.CPU_Dmem_value_a5[4][10] ;
 wire \core.CPU_Dmem_value_a5[4][11] ;
 wire \core.CPU_Dmem_value_a5[4][12] ;
 wire \core.CPU_Dmem_value_a5[4][13] ;
 wire \core.CPU_Dmem_value_a5[4][14] ;
 wire \core.CPU_Dmem_value_a5[4][15] ;
 wire \core.CPU_Dmem_value_a5[4][16] ;
 wire \core.CPU_Dmem_value_a5[4][17] ;
 wire \core.CPU_Dmem_value_a5[4][18] ;
 wire \core.CPU_Dmem_value_a5[4][19] ;
 wire \core.CPU_Dmem_value_a5[4][1] ;
 wire \core.CPU_Dmem_value_a5[4][20] ;
 wire \core.CPU_Dmem_value_a5[4][21] ;
 wire \core.CPU_Dmem_value_a5[4][22] ;
 wire \core.CPU_Dmem_value_a5[4][23] ;
 wire \core.CPU_Dmem_value_a5[4][24] ;
 wire \core.CPU_Dmem_value_a5[4][25] ;
 wire \core.CPU_Dmem_value_a5[4][26] ;
 wire \core.CPU_Dmem_value_a5[4][27] ;
 wire \core.CPU_Dmem_value_a5[4][28] ;
 wire \core.CPU_Dmem_value_a5[4][29] ;
 wire \core.CPU_Dmem_value_a5[4][2] ;
 wire \core.CPU_Dmem_value_a5[4][30] ;
 wire \core.CPU_Dmem_value_a5[4][31] ;
 wire \core.CPU_Dmem_value_a5[4][3] ;
 wire \core.CPU_Dmem_value_a5[4][4] ;
 wire \core.CPU_Dmem_value_a5[4][5] ;
 wire \core.CPU_Dmem_value_a5[4][6] ;
 wire \core.CPU_Dmem_value_a5[4][7] ;
 wire \core.CPU_Dmem_value_a5[4][8] ;
 wire \core.CPU_Dmem_value_a5[4][9] ;
 wire \core.CPU_Dmem_value_a5[5][0] ;
 wire \core.CPU_Dmem_value_a5[5][10] ;
 wire \core.CPU_Dmem_value_a5[5][11] ;
 wire \core.CPU_Dmem_value_a5[5][12] ;
 wire \core.CPU_Dmem_value_a5[5][13] ;
 wire \core.CPU_Dmem_value_a5[5][14] ;
 wire \core.CPU_Dmem_value_a5[5][15] ;
 wire \core.CPU_Dmem_value_a5[5][16] ;
 wire \core.CPU_Dmem_value_a5[5][17] ;
 wire \core.CPU_Dmem_value_a5[5][18] ;
 wire \core.CPU_Dmem_value_a5[5][19] ;
 wire \core.CPU_Dmem_value_a5[5][1] ;
 wire \core.CPU_Dmem_value_a5[5][20] ;
 wire \core.CPU_Dmem_value_a5[5][21] ;
 wire \core.CPU_Dmem_value_a5[5][22] ;
 wire \core.CPU_Dmem_value_a5[5][23] ;
 wire \core.CPU_Dmem_value_a5[5][24] ;
 wire \core.CPU_Dmem_value_a5[5][25] ;
 wire \core.CPU_Dmem_value_a5[5][26] ;
 wire \core.CPU_Dmem_value_a5[5][27] ;
 wire \core.CPU_Dmem_value_a5[5][28] ;
 wire \core.CPU_Dmem_value_a5[5][29] ;
 wire \core.CPU_Dmem_value_a5[5][2] ;
 wire \core.CPU_Dmem_value_a5[5][30] ;
 wire \core.CPU_Dmem_value_a5[5][31] ;
 wire \core.CPU_Dmem_value_a5[5][3] ;
 wire \core.CPU_Dmem_value_a5[5][4] ;
 wire \core.CPU_Dmem_value_a5[5][5] ;
 wire \core.CPU_Dmem_value_a5[5][6] ;
 wire \core.CPU_Dmem_value_a5[5][7] ;
 wire \core.CPU_Dmem_value_a5[5][8] ;
 wire \core.CPU_Dmem_value_a5[5][9] ;
 wire \core.CPU_Dmem_value_a5[6][0] ;
 wire \core.CPU_Dmem_value_a5[6][10] ;
 wire \core.CPU_Dmem_value_a5[6][11] ;
 wire \core.CPU_Dmem_value_a5[6][12] ;
 wire \core.CPU_Dmem_value_a5[6][13] ;
 wire \core.CPU_Dmem_value_a5[6][14] ;
 wire \core.CPU_Dmem_value_a5[6][15] ;
 wire \core.CPU_Dmem_value_a5[6][16] ;
 wire \core.CPU_Dmem_value_a5[6][17] ;
 wire \core.CPU_Dmem_value_a5[6][18] ;
 wire \core.CPU_Dmem_value_a5[6][19] ;
 wire \core.CPU_Dmem_value_a5[6][1] ;
 wire \core.CPU_Dmem_value_a5[6][20] ;
 wire \core.CPU_Dmem_value_a5[6][21] ;
 wire \core.CPU_Dmem_value_a5[6][22] ;
 wire \core.CPU_Dmem_value_a5[6][23] ;
 wire \core.CPU_Dmem_value_a5[6][24] ;
 wire \core.CPU_Dmem_value_a5[6][25] ;
 wire \core.CPU_Dmem_value_a5[6][26] ;
 wire \core.CPU_Dmem_value_a5[6][27] ;
 wire \core.CPU_Dmem_value_a5[6][28] ;
 wire \core.CPU_Dmem_value_a5[6][29] ;
 wire \core.CPU_Dmem_value_a5[6][2] ;
 wire \core.CPU_Dmem_value_a5[6][30] ;
 wire \core.CPU_Dmem_value_a5[6][31] ;
 wire \core.CPU_Dmem_value_a5[6][3] ;
 wire \core.CPU_Dmem_value_a5[6][4] ;
 wire \core.CPU_Dmem_value_a5[6][5] ;
 wire \core.CPU_Dmem_value_a5[6][6] ;
 wire \core.CPU_Dmem_value_a5[6][7] ;
 wire \core.CPU_Dmem_value_a5[6][8] ;
 wire \core.CPU_Dmem_value_a5[6][9] ;
 wire \core.CPU_Dmem_value_a5[7][0] ;
 wire \core.CPU_Dmem_value_a5[7][10] ;
 wire \core.CPU_Dmem_value_a5[7][11] ;
 wire \core.CPU_Dmem_value_a5[7][12] ;
 wire \core.CPU_Dmem_value_a5[7][13] ;
 wire \core.CPU_Dmem_value_a5[7][14] ;
 wire \core.CPU_Dmem_value_a5[7][15] ;
 wire \core.CPU_Dmem_value_a5[7][16] ;
 wire \core.CPU_Dmem_value_a5[7][17] ;
 wire \core.CPU_Dmem_value_a5[7][18] ;
 wire \core.CPU_Dmem_value_a5[7][19] ;
 wire \core.CPU_Dmem_value_a5[7][1] ;
 wire \core.CPU_Dmem_value_a5[7][20] ;
 wire \core.CPU_Dmem_value_a5[7][21] ;
 wire \core.CPU_Dmem_value_a5[7][22] ;
 wire \core.CPU_Dmem_value_a5[7][23] ;
 wire \core.CPU_Dmem_value_a5[7][24] ;
 wire \core.CPU_Dmem_value_a5[7][25] ;
 wire \core.CPU_Dmem_value_a5[7][26] ;
 wire \core.CPU_Dmem_value_a5[7][27] ;
 wire \core.CPU_Dmem_value_a5[7][28] ;
 wire \core.CPU_Dmem_value_a5[7][29] ;
 wire \core.CPU_Dmem_value_a5[7][2] ;
 wire \core.CPU_Dmem_value_a5[7][30] ;
 wire \core.CPU_Dmem_value_a5[7][31] ;
 wire \core.CPU_Dmem_value_a5[7][3] ;
 wire \core.CPU_Dmem_value_a5[7][4] ;
 wire \core.CPU_Dmem_value_a5[7][5] ;
 wire \core.CPU_Dmem_value_a5[7][6] ;
 wire \core.CPU_Dmem_value_a5[7][7] ;
 wire \core.CPU_Dmem_value_a5[7][8] ;
 wire \core.CPU_Dmem_value_a5[7][9] ;
 wire \core.CPU_Dmem_value_a5[8][0] ;
 wire \core.CPU_Dmem_value_a5[8][10] ;
 wire \core.CPU_Dmem_value_a5[8][11] ;
 wire \core.CPU_Dmem_value_a5[8][12] ;
 wire \core.CPU_Dmem_value_a5[8][13] ;
 wire \core.CPU_Dmem_value_a5[8][14] ;
 wire \core.CPU_Dmem_value_a5[8][15] ;
 wire \core.CPU_Dmem_value_a5[8][16] ;
 wire \core.CPU_Dmem_value_a5[8][17] ;
 wire \core.CPU_Dmem_value_a5[8][18] ;
 wire \core.CPU_Dmem_value_a5[8][19] ;
 wire \core.CPU_Dmem_value_a5[8][1] ;
 wire \core.CPU_Dmem_value_a5[8][20] ;
 wire \core.CPU_Dmem_value_a5[8][21] ;
 wire \core.CPU_Dmem_value_a5[8][22] ;
 wire \core.CPU_Dmem_value_a5[8][23] ;
 wire \core.CPU_Dmem_value_a5[8][24] ;
 wire \core.CPU_Dmem_value_a5[8][25] ;
 wire \core.CPU_Dmem_value_a5[8][26] ;
 wire \core.CPU_Dmem_value_a5[8][27] ;
 wire \core.CPU_Dmem_value_a5[8][28] ;
 wire \core.CPU_Dmem_value_a5[8][29] ;
 wire \core.CPU_Dmem_value_a5[8][2] ;
 wire \core.CPU_Dmem_value_a5[8][30] ;
 wire \core.CPU_Dmem_value_a5[8][31] ;
 wire \core.CPU_Dmem_value_a5[8][3] ;
 wire \core.CPU_Dmem_value_a5[8][4] ;
 wire \core.CPU_Dmem_value_a5[8][5] ;
 wire \core.CPU_Dmem_value_a5[8][6] ;
 wire \core.CPU_Dmem_value_a5[8][7] ;
 wire \core.CPU_Dmem_value_a5[8][8] ;
 wire \core.CPU_Dmem_value_a5[8][9] ;
 wire \core.CPU_Dmem_value_a5[9][0] ;
 wire \core.CPU_Dmem_value_a5[9][10] ;
 wire \core.CPU_Dmem_value_a5[9][11] ;
 wire \core.CPU_Dmem_value_a5[9][12] ;
 wire \core.CPU_Dmem_value_a5[9][13] ;
 wire \core.CPU_Dmem_value_a5[9][14] ;
 wire \core.CPU_Dmem_value_a5[9][15] ;
 wire \core.CPU_Dmem_value_a5[9][16] ;
 wire \core.CPU_Dmem_value_a5[9][17] ;
 wire \core.CPU_Dmem_value_a5[9][18] ;
 wire \core.CPU_Dmem_value_a5[9][19] ;
 wire \core.CPU_Dmem_value_a5[9][1] ;
 wire \core.CPU_Dmem_value_a5[9][20] ;
 wire \core.CPU_Dmem_value_a5[9][21] ;
 wire \core.CPU_Dmem_value_a5[9][22] ;
 wire \core.CPU_Dmem_value_a5[9][23] ;
 wire \core.CPU_Dmem_value_a5[9][24] ;
 wire \core.CPU_Dmem_value_a5[9][25] ;
 wire \core.CPU_Dmem_value_a5[9][26] ;
 wire \core.CPU_Dmem_value_a5[9][27] ;
 wire \core.CPU_Dmem_value_a5[9][28] ;
 wire \core.CPU_Dmem_value_a5[9][29] ;
 wire \core.CPU_Dmem_value_a5[9][2] ;
 wire \core.CPU_Dmem_value_a5[9][30] ;
 wire \core.CPU_Dmem_value_a5[9][31] ;
 wire \core.CPU_Dmem_value_a5[9][3] ;
 wire \core.CPU_Dmem_value_a5[9][4] ;
 wire \core.CPU_Dmem_value_a5[9][5] ;
 wire \core.CPU_Dmem_value_a5[9][6] ;
 wire \core.CPU_Dmem_value_a5[9][7] ;
 wire \core.CPU_Dmem_value_a5[9][8] ;
 wire \core.CPU_Dmem_value_a5[9][9] ;
 wire \core.CPU_Xreg_value_a4[0][0] ;
 wire \core.CPU_Xreg_value_a4[0][10] ;
 wire \core.CPU_Xreg_value_a4[0][11] ;
 wire \core.CPU_Xreg_value_a4[0][12] ;
 wire \core.CPU_Xreg_value_a4[0][13] ;
 wire \core.CPU_Xreg_value_a4[0][14] ;
 wire \core.CPU_Xreg_value_a4[0][15] ;
 wire \core.CPU_Xreg_value_a4[0][16] ;
 wire \core.CPU_Xreg_value_a4[0][17] ;
 wire \core.CPU_Xreg_value_a4[0][18] ;
 wire \core.CPU_Xreg_value_a4[0][19] ;
 wire \core.CPU_Xreg_value_a4[0][1] ;
 wire \core.CPU_Xreg_value_a4[0][20] ;
 wire \core.CPU_Xreg_value_a4[0][21] ;
 wire \core.CPU_Xreg_value_a4[0][22] ;
 wire \core.CPU_Xreg_value_a4[0][23] ;
 wire \core.CPU_Xreg_value_a4[0][24] ;
 wire \core.CPU_Xreg_value_a4[0][25] ;
 wire \core.CPU_Xreg_value_a4[0][26] ;
 wire \core.CPU_Xreg_value_a4[0][27] ;
 wire \core.CPU_Xreg_value_a4[0][28] ;
 wire \core.CPU_Xreg_value_a4[0][29] ;
 wire \core.CPU_Xreg_value_a4[0][2] ;
 wire \core.CPU_Xreg_value_a4[0][30] ;
 wire \core.CPU_Xreg_value_a4[0][31] ;
 wire \core.CPU_Xreg_value_a4[0][3] ;
 wire \core.CPU_Xreg_value_a4[0][4] ;
 wire \core.CPU_Xreg_value_a4[0][5] ;
 wire \core.CPU_Xreg_value_a4[0][6] ;
 wire \core.CPU_Xreg_value_a4[0][7] ;
 wire \core.CPU_Xreg_value_a4[0][8] ;
 wire \core.CPU_Xreg_value_a4[0][9] ;
 wire \core.CPU_Xreg_value_a4[10][0] ;
 wire \core.CPU_Xreg_value_a4[10][10] ;
 wire \core.CPU_Xreg_value_a4[10][11] ;
 wire \core.CPU_Xreg_value_a4[10][12] ;
 wire \core.CPU_Xreg_value_a4[10][13] ;
 wire \core.CPU_Xreg_value_a4[10][14] ;
 wire \core.CPU_Xreg_value_a4[10][15] ;
 wire \core.CPU_Xreg_value_a4[10][16] ;
 wire \core.CPU_Xreg_value_a4[10][17] ;
 wire \core.CPU_Xreg_value_a4[10][18] ;
 wire \core.CPU_Xreg_value_a4[10][19] ;
 wire \core.CPU_Xreg_value_a4[10][1] ;
 wire \core.CPU_Xreg_value_a4[10][20] ;
 wire \core.CPU_Xreg_value_a4[10][21] ;
 wire \core.CPU_Xreg_value_a4[10][22] ;
 wire \core.CPU_Xreg_value_a4[10][23] ;
 wire \core.CPU_Xreg_value_a4[10][24] ;
 wire \core.CPU_Xreg_value_a4[10][25] ;
 wire \core.CPU_Xreg_value_a4[10][26] ;
 wire \core.CPU_Xreg_value_a4[10][27] ;
 wire \core.CPU_Xreg_value_a4[10][28] ;
 wire \core.CPU_Xreg_value_a4[10][29] ;
 wire \core.CPU_Xreg_value_a4[10][2] ;
 wire \core.CPU_Xreg_value_a4[10][30] ;
 wire \core.CPU_Xreg_value_a4[10][31] ;
 wire \core.CPU_Xreg_value_a4[10][3] ;
 wire \core.CPU_Xreg_value_a4[10][4] ;
 wire \core.CPU_Xreg_value_a4[10][5] ;
 wire \core.CPU_Xreg_value_a4[10][6] ;
 wire \core.CPU_Xreg_value_a4[10][7] ;
 wire \core.CPU_Xreg_value_a4[10][8] ;
 wire \core.CPU_Xreg_value_a4[10][9] ;
 wire \core.CPU_Xreg_value_a4[11][0] ;
 wire \core.CPU_Xreg_value_a4[11][10] ;
 wire \core.CPU_Xreg_value_a4[11][11] ;
 wire \core.CPU_Xreg_value_a4[11][12] ;
 wire \core.CPU_Xreg_value_a4[11][13] ;
 wire \core.CPU_Xreg_value_a4[11][14] ;
 wire \core.CPU_Xreg_value_a4[11][15] ;
 wire \core.CPU_Xreg_value_a4[11][16] ;
 wire \core.CPU_Xreg_value_a4[11][17] ;
 wire \core.CPU_Xreg_value_a4[11][18] ;
 wire \core.CPU_Xreg_value_a4[11][19] ;
 wire \core.CPU_Xreg_value_a4[11][1] ;
 wire \core.CPU_Xreg_value_a4[11][20] ;
 wire \core.CPU_Xreg_value_a4[11][21] ;
 wire \core.CPU_Xreg_value_a4[11][22] ;
 wire \core.CPU_Xreg_value_a4[11][23] ;
 wire \core.CPU_Xreg_value_a4[11][24] ;
 wire \core.CPU_Xreg_value_a4[11][25] ;
 wire \core.CPU_Xreg_value_a4[11][26] ;
 wire \core.CPU_Xreg_value_a4[11][27] ;
 wire \core.CPU_Xreg_value_a4[11][28] ;
 wire \core.CPU_Xreg_value_a4[11][29] ;
 wire \core.CPU_Xreg_value_a4[11][2] ;
 wire \core.CPU_Xreg_value_a4[11][30] ;
 wire \core.CPU_Xreg_value_a4[11][31] ;
 wire \core.CPU_Xreg_value_a4[11][3] ;
 wire \core.CPU_Xreg_value_a4[11][4] ;
 wire \core.CPU_Xreg_value_a4[11][5] ;
 wire \core.CPU_Xreg_value_a4[11][6] ;
 wire \core.CPU_Xreg_value_a4[11][7] ;
 wire \core.CPU_Xreg_value_a4[11][8] ;
 wire \core.CPU_Xreg_value_a4[11][9] ;
 wire \core.CPU_Xreg_value_a4[16][0] ;
 wire \core.CPU_Xreg_value_a4[16][10] ;
 wire \core.CPU_Xreg_value_a4[16][11] ;
 wire \core.CPU_Xreg_value_a4[16][12] ;
 wire \core.CPU_Xreg_value_a4[16][13] ;
 wire \core.CPU_Xreg_value_a4[16][14] ;
 wire \core.CPU_Xreg_value_a4[16][15] ;
 wire \core.CPU_Xreg_value_a4[16][16] ;
 wire \core.CPU_Xreg_value_a4[16][17] ;
 wire \core.CPU_Xreg_value_a4[16][18] ;
 wire \core.CPU_Xreg_value_a4[16][19] ;
 wire \core.CPU_Xreg_value_a4[16][1] ;
 wire \core.CPU_Xreg_value_a4[16][20] ;
 wire \core.CPU_Xreg_value_a4[16][21] ;
 wire \core.CPU_Xreg_value_a4[16][22] ;
 wire \core.CPU_Xreg_value_a4[16][23] ;
 wire \core.CPU_Xreg_value_a4[16][24] ;
 wire \core.CPU_Xreg_value_a4[16][25] ;
 wire \core.CPU_Xreg_value_a4[16][26] ;
 wire \core.CPU_Xreg_value_a4[16][27] ;
 wire \core.CPU_Xreg_value_a4[16][28] ;
 wire \core.CPU_Xreg_value_a4[16][29] ;
 wire \core.CPU_Xreg_value_a4[16][2] ;
 wire \core.CPU_Xreg_value_a4[16][30] ;
 wire \core.CPU_Xreg_value_a4[16][31] ;
 wire \core.CPU_Xreg_value_a4[16][3] ;
 wire \core.CPU_Xreg_value_a4[16][4] ;
 wire \core.CPU_Xreg_value_a4[16][5] ;
 wire \core.CPU_Xreg_value_a4[16][6] ;
 wire \core.CPU_Xreg_value_a4[16][7] ;
 wire \core.CPU_Xreg_value_a4[16][8] ;
 wire \core.CPU_Xreg_value_a4[16][9] ;
 wire \core.CPU_Xreg_value_a4[17][0] ;
 wire \core.CPU_Xreg_value_a4[17][10] ;
 wire \core.CPU_Xreg_value_a4[17][11] ;
 wire \core.CPU_Xreg_value_a4[17][12] ;
 wire \core.CPU_Xreg_value_a4[17][13] ;
 wire \core.CPU_Xreg_value_a4[17][14] ;
 wire \core.CPU_Xreg_value_a4[17][15] ;
 wire \core.CPU_Xreg_value_a4[17][16] ;
 wire \core.CPU_Xreg_value_a4[17][17] ;
 wire \core.CPU_Xreg_value_a4[17][18] ;
 wire \core.CPU_Xreg_value_a4[17][19] ;
 wire \core.CPU_Xreg_value_a4[17][1] ;
 wire \core.CPU_Xreg_value_a4[17][20] ;
 wire \core.CPU_Xreg_value_a4[17][21] ;
 wire \core.CPU_Xreg_value_a4[17][22] ;
 wire \core.CPU_Xreg_value_a4[17][23] ;
 wire \core.CPU_Xreg_value_a4[17][24] ;
 wire \core.CPU_Xreg_value_a4[17][25] ;
 wire \core.CPU_Xreg_value_a4[17][26] ;
 wire \core.CPU_Xreg_value_a4[17][27] ;
 wire \core.CPU_Xreg_value_a4[17][28] ;
 wire \core.CPU_Xreg_value_a4[17][29] ;
 wire \core.CPU_Xreg_value_a4[17][2] ;
 wire \core.CPU_Xreg_value_a4[17][30] ;
 wire \core.CPU_Xreg_value_a4[17][31] ;
 wire \core.CPU_Xreg_value_a4[17][3] ;
 wire \core.CPU_Xreg_value_a4[17][4] ;
 wire \core.CPU_Xreg_value_a4[17][5] ;
 wire \core.CPU_Xreg_value_a4[17][6] ;
 wire \core.CPU_Xreg_value_a4[17][7] ;
 wire \core.CPU_Xreg_value_a4[17][8] ;
 wire \core.CPU_Xreg_value_a4[17][9] ;
 wire \core.CPU_Xreg_value_a4[1][0] ;
 wire \core.CPU_Xreg_value_a4[1][10] ;
 wire \core.CPU_Xreg_value_a4[1][11] ;
 wire \core.CPU_Xreg_value_a4[1][12] ;
 wire \core.CPU_Xreg_value_a4[1][13] ;
 wire \core.CPU_Xreg_value_a4[1][14] ;
 wire \core.CPU_Xreg_value_a4[1][15] ;
 wire \core.CPU_Xreg_value_a4[1][16] ;
 wire \core.CPU_Xreg_value_a4[1][17] ;
 wire \core.CPU_Xreg_value_a4[1][18] ;
 wire \core.CPU_Xreg_value_a4[1][19] ;
 wire \core.CPU_Xreg_value_a4[1][1] ;
 wire \core.CPU_Xreg_value_a4[1][20] ;
 wire \core.CPU_Xreg_value_a4[1][21] ;
 wire \core.CPU_Xreg_value_a4[1][22] ;
 wire \core.CPU_Xreg_value_a4[1][23] ;
 wire \core.CPU_Xreg_value_a4[1][24] ;
 wire \core.CPU_Xreg_value_a4[1][25] ;
 wire \core.CPU_Xreg_value_a4[1][26] ;
 wire \core.CPU_Xreg_value_a4[1][27] ;
 wire \core.CPU_Xreg_value_a4[1][28] ;
 wire \core.CPU_Xreg_value_a4[1][29] ;
 wire \core.CPU_Xreg_value_a4[1][2] ;
 wire \core.CPU_Xreg_value_a4[1][30] ;
 wire \core.CPU_Xreg_value_a4[1][31] ;
 wire \core.CPU_Xreg_value_a4[1][3] ;
 wire \core.CPU_Xreg_value_a4[1][4] ;
 wire \core.CPU_Xreg_value_a4[1][5] ;
 wire \core.CPU_Xreg_value_a4[1][6] ;
 wire \core.CPU_Xreg_value_a4[1][7] ;
 wire \core.CPU_Xreg_value_a4[1][8] ;
 wire \core.CPU_Xreg_value_a4[1][9] ;
 wire \core.CPU_Xreg_value_a4[26][0] ;
 wire \core.CPU_Xreg_value_a4[26][10] ;
 wire \core.CPU_Xreg_value_a4[26][11] ;
 wire \core.CPU_Xreg_value_a4[26][12] ;
 wire \core.CPU_Xreg_value_a4[26][13] ;
 wire \core.CPU_Xreg_value_a4[26][14] ;
 wire \core.CPU_Xreg_value_a4[26][15] ;
 wire \core.CPU_Xreg_value_a4[26][16] ;
 wire \core.CPU_Xreg_value_a4[26][17] ;
 wire \core.CPU_Xreg_value_a4[26][18] ;
 wire \core.CPU_Xreg_value_a4[26][19] ;
 wire \core.CPU_Xreg_value_a4[26][1] ;
 wire \core.CPU_Xreg_value_a4[26][20] ;
 wire \core.CPU_Xreg_value_a4[26][21] ;
 wire \core.CPU_Xreg_value_a4[26][22] ;
 wire \core.CPU_Xreg_value_a4[26][23] ;
 wire \core.CPU_Xreg_value_a4[26][24] ;
 wire \core.CPU_Xreg_value_a4[26][25] ;
 wire \core.CPU_Xreg_value_a4[26][26] ;
 wire \core.CPU_Xreg_value_a4[26][27] ;
 wire \core.CPU_Xreg_value_a4[26][28] ;
 wire \core.CPU_Xreg_value_a4[26][29] ;
 wire \core.CPU_Xreg_value_a4[26][2] ;
 wire \core.CPU_Xreg_value_a4[26][30] ;
 wire \core.CPU_Xreg_value_a4[26][31] ;
 wire \core.CPU_Xreg_value_a4[26][3] ;
 wire \core.CPU_Xreg_value_a4[26][4] ;
 wire \core.CPU_Xreg_value_a4[26][5] ;
 wire \core.CPU_Xreg_value_a4[26][6] ;
 wire \core.CPU_Xreg_value_a4[26][7] ;
 wire \core.CPU_Xreg_value_a4[26][8] ;
 wire \core.CPU_Xreg_value_a4[26][9] ;
 wire \core.CPU_Xreg_value_a4[27][0] ;
 wire \core.CPU_Xreg_value_a4[27][10] ;
 wire \core.CPU_Xreg_value_a4[27][11] ;
 wire \core.CPU_Xreg_value_a4[27][12] ;
 wire \core.CPU_Xreg_value_a4[27][13] ;
 wire \core.CPU_Xreg_value_a4[27][14] ;
 wire \core.CPU_Xreg_value_a4[27][15] ;
 wire \core.CPU_Xreg_value_a4[27][16] ;
 wire \core.CPU_Xreg_value_a4[27][17] ;
 wire \core.CPU_Xreg_value_a4[27][18] ;
 wire \core.CPU_Xreg_value_a4[27][19] ;
 wire \core.CPU_Xreg_value_a4[27][1] ;
 wire \core.CPU_Xreg_value_a4[27][20] ;
 wire \core.CPU_Xreg_value_a4[27][21] ;
 wire \core.CPU_Xreg_value_a4[27][22] ;
 wire \core.CPU_Xreg_value_a4[27][23] ;
 wire \core.CPU_Xreg_value_a4[27][24] ;
 wire \core.CPU_Xreg_value_a4[27][25] ;
 wire \core.CPU_Xreg_value_a4[27][26] ;
 wire \core.CPU_Xreg_value_a4[27][27] ;
 wire \core.CPU_Xreg_value_a4[27][28] ;
 wire \core.CPU_Xreg_value_a4[27][29] ;
 wire \core.CPU_Xreg_value_a4[27][2] ;
 wire \core.CPU_Xreg_value_a4[27][30] ;
 wire \core.CPU_Xreg_value_a4[27][31] ;
 wire \core.CPU_Xreg_value_a4[27][3] ;
 wire \core.CPU_Xreg_value_a4[27][4] ;
 wire \core.CPU_Xreg_value_a4[27][5] ;
 wire \core.CPU_Xreg_value_a4[27][6] ;
 wire \core.CPU_Xreg_value_a4[27][7] ;
 wire \core.CPU_Xreg_value_a4[27][8] ;
 wire \core.CPU_Xreg_value_a4[27][9] ;
 wire \core.CPU_Xreg_value_a4[2][0] ;
 wire \core.CPU_Xreg_value_a4[2][10] ;
 wire \core.CPU_Xreg_value_a4[2][11] ;
 wire \core.CPU_Xreg_value_a4[2][12] ;
 wire \core.CPU_Xreg_value_a4[2][13] ;
 wire \core.CPU_Xreg_value_a4[2][14] ;
 wire \core.CPU_Xreg_value_a4[2][15] ;
 wire \core.CPU_Xreg_value_a4[2][16] ;
 wire \core.CPU_Xreg_value_a4[2][17] ;
 wire \core.CPU_Xreg_value_a4[2][18] ;
 wire \core.CPU_Xreg_value_a4[2][19] ;
 wire \core.CPU_Xreg_value_a4[2][1] ;
 wire \core.CPU_Xreg_value_a4[2][20] ;
 wire \core.CPU_Xreg_value_a4[2][21] ;
 wire \core.CPU_Xreg_value_a4[2][22] ;
 wire \core.CPU_Xreg_value_a4[2][23] ;
 wire \core.CPU_Xreg_value_a4[2][24] ;
 wire \core.CPU_Xreg_value_a4[2][25] ;
 wire \core.CPU_Xreg_value_a4[2][26] ;
 wire \core.CPU_Xreg_value_a4[2][27] ;
 wire \core.CPU_Xreg_value_a4[2][28] ;
 wire \core.CPU_Xreg_value_a4[2][29] ;
 wire \core.CPU_Xreg_value_a4[2][2] ;
 wire \core.CPU_Xreg_value_a4[2][30] ;
 wire \core.CPU_Xreg_value_a4[2][31] ;
 wire \core.CPU_Xreg_value_a4[2][3] ;
 wire \core.CPU_Xreg_value_a4[2][4] ;
 wire \core.CPU_Xreg_value_a4[2][5] ;
 wire \core.CPU_Xreg_value_a4[2][6] ;
 wire \core.CPU_Xreg_value_a4[2][7] ;
 wire \core.CPU_Xreg_value_a4[2][8] ;
 wire \core.CPU_Xreg_value_a4[2][9] ;
 wire \core.CPU_Xreg_value_a4[3][0] ;
 wire \core.CPU_Xreg_value_a4[3][10] ;
 wire \core.CPU_Xreg_value_a4[3][11] ;
 wire \core.CPU_Xreg_value_a4[3][12] ;
 wire \core.CPU_Xreg_value_a4[3][13] ;
 wire \core.CPU_Xreg_value_a4[3][14] ;
 wire \core.CPU_Xreg_value_a4[3][15] ;
 wire \core.CPU_Xreg_value_a4[3][16] ;
 wire \core.CPU_Xreg_value_a4[3][17] ;
 wire \core.CPU_Xreg_value_a4[3][18] ;
 wire \core.CPU_Xreg_value_a4[3][19] ;
 wire \core.CPU_Xreg_value_a4[3][1] ;
 wire \core.CPU_Xreg_value_a4[3][20] ;
 wire \core.CPU_Xreg_value_a4[3][21] ;
 wire \core.CPU_Xreg_value_a4[3][22] ;
 wire \core.CPU_Xreg_value_a4[3][23] ;
 wire \core.CPU_Xreg_value_a4[3][24] ;
 wire \core.CPU_Xreg_value_a4[3][25] ;
 wire \core.CPU_Xreg_value_a4[3][26] ;
 wire \core.CPU_Xreg_value_a4[3][27] ;
 wire \core.CPU_Xreg_value_a4[3][28] ;
 wire \core.CPU_Xreg_value_a4[3][29] ;
 wire \core.CPU_Xreg_value_a4[3][2] ;
 wire \core.CPU_Xreg_value_a4[3][30] ;
 wire \core.CPU_Xreg_value_a4[3][31] ;
 wire \core.CPU_Xreg_value_a4[3][3] ;
 wire \core.CPU_Xreg_value_a4[3][4] ;
 wire \core.CPU_Xreg_value_a4[3][5] ;
 wire \core.CPU_Xreg_value_a4[3][6] ;
 wire \core.CPU_Xreg_value_a4[3][7] ;
 wire \core.CPU_Xreg_value_a4[3][8] ;
 wire \core.CPU_Xreg_value_a4[3][9] ;
 wire \core.CPU_Xreg_value_a4[8][0] ;
 wire \core.CPU_Xreg_value_a4[8][10] ;
 wire \core.CPU_Xreg_value_a4[8][11] ;
 wire \core.CPU_Xreg_value_a4[8][12] ;
 wire \core.CPU_Xreg_value_a4[8][13] ;
 wire \core.CPU_Xreg_value_a4[8][14] ;
 wire \core.CPU_Xreg_value_a4[8][15] ;
 wire \core.CPU_Xreg_value_a4[8][16] ;
 wire \core.CPU_Xreg_value_a4[8][17] ;
 wire \core.CPU_Xreg_value_a4[8][18] ;
 wire \core.CPU_Xreg_value_a4[8][19] ;
 wire \core.CPU_Xreg_value_a4[8][1] ;
 wire \core.CPU_Xreg_value_a4[8][20] ;
 wire \core.CPU_Xreg_value_a4[8][21] ;
 wire \core.CPU_Xreg_value_a4[8][22] ;
 wire \core.CPU_Xreg_value_a4[8][23] ;
 wire \core.CPU_Xreg_value_a4[8][24] ;
 wire \core.CPU_Xreg_value_a4[8][25] ;
 wire \core.CPU_Xreg_value_a4[8][26] ;
 wire \core.CPU_Xreg_value_a4[8][27] ;
 wire \core.CPU_Xreg_value_a4[8][28] ;
 wire \core.CPU_Xreg_value_a4[8][29] ;
 wire \core.CPU_Xreg_value_a4[8][2] ;
 wire \core.CPU_Xreg_value_a4[8][30] ;
 wire \core.CPU_Xreg_value_a4[8][31] ;
 wire \core.CPU_Xreg_value_a4[8][3] ;
 wire \core.CPU_Xreg_value_a4[8][4] ;
 wire \core.CPU_Xreg_value_a4[8][5] ;
 wire \core.CPU_Xreg_value_a4[8][6] ;
 wire \core.CPU_Xreg_value_a4[8][7] ;
 wire \core.CPU_Xreg_value_a4[8][8] ;
 wire \core.CPU_Xreg_value_a4[8][9] ;
 wire \core.CPU_Xreg_value_a4[9][0] ;
 wire \core.CPU_Xreg_value_a4[9][10] ;
 wire \core.CPU_Xreg_value_a4[9][11] ;
 wire \core.CPU_Xreg_value_a4[9][12] ;
 wire \core.CPU_Xreg_value_a4[9][13] ;
 wire \core.CPU_Xreg_value_a4[9][14] ;
 wire \core.CPU_Xreg_value_a4[9][15] ;
 wire \core.CPU_Xreg_value_a4[9][16] ;
 wire \core.CPU_Xreg_value_a4[9][17] ;
 wire \core.CPU_Xreg_value_a4[9][18] ;
 wire \core.CPU_Xreg_value_a4[9][19] ;
 wire \core.CPU_Xreg_value_a4[9][1] ;
 wire \core.CPU_Xreg_value_a4[9][20] ;
 wire \core.CPU_Xreg_value_a4[9][21] ;
 wire \core.CPU_Xreg_value_a4[9][22] ;
 wire \core.CPU_Xreg_value_a4[9][23] ;
 wire \core.CPU_Xreg_value_a4[9][24] ;
 wire \core.CPU_Xreg_value_a4[9][25] ;
 wire \core.CPU_Xreg_value_a4[9][26] ;
 wire \core.CPU_Xreg_value_a4[9][27] ;
 wire \core.CPU_Xreg_value_a4[9][28] ;
 wire \core.CPU_Xreg_value_a4[9][29] ;
 wire \core.CPU_Xreg_value_a4[9][2] ;
 wire \core.CPU_Xreg_value_a4[9][30] ;
 wire \core.CPU_Xreg_value_a4[9][31] ;
 wire \core.CPU_Xreg_value_a4[9][3] ;
 wire \core.CPU_Xreg_value_a4[9][4] ;
 wire \core.CPU_Xreg_value_a4[9][5] ;
 wire \core.CPU_Xreg_value_a4[9][6] ;
 wire \core.CPU_Xreg_value_a4[9][7] ;
 wire \core.CPU_Xreg_value_a4[9][8] ;
 wire \core.CPU_Xreg_value_a4[9][9] ;
 wire \core.CPU_Xreg_value_a5[17][0] ;
 wire \core.CPU_Xreg_value_a5[17][1] ;
 wire \core.CPU_Xreg_value_a5[17][2] ;
 wire \core.CPU_Xreg_value_a5[17][3] ;
 wire \core.CPU_Xreg_value_a5[17][4] ;
 wire \core.CPU_Xreg_value_a5[17][5] ;
 wire \core.CPU_Xreg_value_a5[17][6] ;
 wire \core.CPU_Xreg_value_a5[17][7] ;
 wire \core.CPU_Xreg_value_a5[17][8] ;
 wire \core.CPU_Xreg_value_a5[17][9] ;
 wire \core.CPU_br_tgt_pc_a2[0] ;
 wire \core.CPU_br_tgt_pc_a2[1] ;
 wire \core.CPU_br_tgt_pc_a2[2] ;
 wire \core.CPU_br_tgt_pc_a2[3] ;
 wire \core.CPU_br_tgt_pc_a2[4] ;
 wire \core.CPU_br_tgt_pc_a2[5] ;
 wire \core.CPU_br_tgt_pc_a3[0] ;
 wire \core.CPU_br_tgt_pc_a3[1] ;
 wire \core.CPU_br_tgt_pc_a3[2] ;
 wire \core.CPU_br_tgt_pc_a3[3] ;
 wire \core.CPU_br_tgt_pc_a3[4] ;
 wire \core.CPU_br_tgt_pc_a3[5] ;
 wire \core.CPU_dmem_addr_a4[0] ;
 wire \core.CPU_dmem_addr_a4[1] ;
 wire \core.CPU_dmem_addr_a4[2] ;
 wire \core.CPU_dmem_addr_a4[3] ;
 wire \core.CPU_dmem_rd_data_a5[0] ;
 wire \core.CPU_dmem_rd_data_a5[10] ;
 wire \core.CPU_dmem_rd_data_a5[11] ;
 wire \core.CPU_dmem_rd_data_a5[12] ;
 wire \core.CPU_dmem_rd_data_a5[13] ;
 wire \core.CPU_dmem_rd_data_a5[14] ;
 wire \core.CPU_dmem_rd_data_a5[15] ;
 wire \core.CPU_dmem_rd_data_a5[16] ;
 wire \core.CPU_dmem_rd_data_a5[17] ;
 wire \core.CPU_dmem_rd_data_a5[18] ;
 wire \core.CPU_dmem_rd_data_a5[19] ;
 wire \core.CPU_dmem_rd_data_a5[1] ;
 wire \core.CPU_dmem_rd_data_a5[20] ;
 wire \core.CPU_dmem_rd_data_a5[21] ;
 wire \core.CPU_dmem_rd_data_a5[22] ;
 wire \core.CPU_dmem_rd_data_a5[23] ;
 wire \core.CPU_dmem_rd_data_a5[24] ;
 wire \core.CPU_dmem_rd_data_a5[25] ;
 wire \core.CPU_dmem_rd_data_a5[26] ;
 wire \core.CPU_dmem_rd_data_a5[27] ;
 wire \core.CPU_dmem_rd_data_a5[28] ;
 wire \core.CPU_dmem_rd_data_a5[29] ;
 wire \core.CPU_dmem_rd_data_a5[2] ;
 wire \core.CPU_dmem_rd_data_a5[30] ;
 wire \core.CPU_dmem_rd_data_a5[31] ;
 wire \core.CPU_dmem_rd_data_a5[3] ;
 wire \core.CPU_dmem_rd_data_a5[4] ;
 wire \core.CPU_dmem_rd_data_a5[5] ;
 wire \core.CPU_dmem_rd_data_a5[6] ;
 wire \core.CPU_dmem_rd_data_a5[7] ;
 wire \core.CPU_dmem_rd_data_a5[8] ;
 wire \core.CPU_dmem_rd_data_a5[9] ;
 wire \core.CPU_dmem_rd_en_a4 ;
 wire \core.CPU_dmem_wr_data_a4[0] ;
 wire \core.CPU_dmem_wr_data_a4[10] ;
 wire \core.CPU_dmem_wr_data_a4[11] ;
 wire \core.CPU_dmem_wr_data_a4[12] ;
 wire \core.CPU_dmem_wr_data_a4[13] ;
 wire \core.CPU_dmem_wr_data_a4[14] ;
 wire \core.CPU_dmem_wr_data_a4[15] ;
 wire \core.CPU_dmem_wr_data_a4[16] ;
 wire \core.CPU_dmem_wr_data_a4[17] ;
 wire \core.CPU_dmem_wr_data_a4[18] ;
 wire \core.CPU_dmem_wr_data_a4[19] ;
 wire \core.CPU_dmem_wr_data_a4[1] ;
 wire \core.CPU_dmem_wr_data_a4[20] ;
 wire \core.CPU_dmem_wr_data_a4[21] ;
 wire \core.CPU_dmem_wr_data_a4[22] ;
 wire \core.CPU_dmem_wr_data_a4[23] ;
 wire \core.CPU_dmem_wr_data_a4[24] ;
 wire \core.CPU_dmem_wr_data_a4[25] ;
 wire \core.CPU_dmem_wr_data_a4[26] ;
 wire \core.CPU_dmem_wr_data_a4[27] ;
 wire \core.CPU_dmem_wr_data_a4[28] ;
 wire \core.CPU_dmem_wr_data_a4[29] ;
 wire \core.CPU_dmem_wr_data_a4[2] ;
 wire \core.CPU_dmem_wr_data_a4[30] ;
 wire \core.CPU_dmem_wr_data_a4[31] ;
 wire \core.CPU_dmem_wr_data_a4[3] ;
 wire \core.CPU_dmem_wr_data_a4[4] ;
 wire \core.CPU_dmem_wr_data_a4[5] ;
 wire \core.CPU_dmem_wr_data_a4[6] ;
 wire \core.CPU_dmem_wr_data_a4[7] ;
 wire \core.CPU_dmem_wr_data_a4[8] ;
 wire \core.CPU_dmem_wr_data_a4[9] ;
 wire \core.CPU_imem_rd_addr_a1[0] ;
 wire \core.CPU_imem_rd_addr_a1[1] ;
 wire \core.CPU_imem_rd_addr_a1[2] ;
 wire \core.CPU_imem_rd_addr_a1[3] ;
 wire \core.CPU_imem_rd_data_a1[10] ;
 wire \core.CPU_imem_rd_data_a1[11] ;
 wire \core.CPU_imem_rd_data_a1[20] ;
 wire \core.CPU_imem_rd_data_a1[21] ;
 wire \core.CPU_imem_rd_data_a1[23] ;
 wire \core.CPU_imem_rd_data_a1[7] ;
 wire \core.CPU_imem_rd_data_a1[8] ;
 wire \core.CPU_imm_a1[0] ;
 wire \core.CPU_imm_a1[10] ;
 wire \core.CPU_imm_a1[11] ;
 wire \core.CPU_imm_a1[12] ;
 wire \core.CPU_imm_a1[1] ;
 wire \core.CPU_imm_a1[3] ;
 wire \core.CPU_imm_a1[5] ;
 wire \core.CPU_imm_a2[0] ;
 wire \core.CPU_imm_a2[10] ;
 wire \core.CPU_imm_a2[11] ;
 wire \core.CPU_imm_a2[12] ;
 wire \core.CPU_imm_a2[1] ;
 wire \core.CPU_imm_a2[3] ;
 wire \core.CPU_imm_a2[4] ;
 wire \core.CPU_imm_a2[5] ;
 wire \core.CPU_imm_a3[0] ;
 wire \core.CPU_imm_a3[10] ;
 wire \core.CPU_imm_a3[11] ;
 wire \core.CPU_imm_a3[12] ;
 wire \core.CPU_imm_a3[1] ;
 wire \core.CPU_imm_a3[3] ;
 wire \core.CPU_imm_a3[4] ;
 wire \core.CPU_imm_a3[5] ;
 wire \core.CPU_inc_pc_a1[0] ;
 wire \core.CPU_inc_pc_a1[1] ;
 wire \core.CPU_inc_pc_a1[2] ;
 wire \core.CPU_inc_pc_a1[3] ;
 wire \core.CPU_inc_pc_a1[4] ;
 wire \core.CPU_inc_pc_a1[5] ;
 wire \core.CPU_inc_pc_a2[0] ;
 wire \core.CPU_inc_pc_a2[1] ;
 wire \core.CPU_inc_pc_a2[2] ;
 wire \core.CPU_inc_pc_a2[3] ;
 wire \core.CPU_inc_pc_a2[4] ;
 wire \core.CPU_inc_pc_a2[5] ;
 wire \core.CPU_inc_pc_a3[0] ;
 wire \core.CPU_inc_pc_a3[1] ;
 wire \core.CPU_inc_pc_a3[2] ;
 wire \core.CPU_inc_pc_a3[3] ;
 wire \core.CPU_inc_pc_a3[4] ;
 wire \core.CPU_inc_pc_a3[5] ;
 wire \core.CPU_is_add_a1 ;
 wire \core.CPU_is_add_a2 ;
 wire \core.CPU_is_add_a3 ;
 wire \core.CPU_is_addi_a1 ;
 wire \core.CPU_is_addi_a2 ;
 wire \core.CPU_is_addi_a3 ;
 wire \core.CPU_is_beq_a1 ;
 wire \core.CPU_is_beq_a2 ;
 wire \core.CPU_is_beq_a3 ;
 wire \core.CPU_is_bne_a1 ;
 wire \core.CPU_is_bne_a2 ;
 wire \core.CPU_is_bne_a3 ;
 wire \core.CPU_is_load_a2 ;
 wire \core.CPU_is_load_a3 ;
 wire \core.CPU_is_s_instr_a2 ;
 wire \core.CPU_is_s_instr_a3 ;
 wire \core.CPU_is_s_instr_a4 ;
 wire \core.CPU_is_sll_a2 ;
 wire \core.CPU_is_sll_a3 ;
 wire \core.CPU_is_slli_a2 ;
 wire \core.CPU_is_slli_a3 ;
 wire \core.CPU_is_sub_a1 ;
 wire \core.CPU_is_sub_a2 ;
 wire \core.CPU_is_sub_a3 ;
 wire \core.CPU_pc_a2[2] ;
 wire \core.CPU_pc_a2[3] ;
 wire \core.CPU_pc_a2[4] ;
 wire \core.CPU_pc_a2[5] ;
 wire \core.CPU_rd_a2[0] ;
 wire \core.CPU_rd_a2[1] ;
 wire \core.CPU_rd_a2[3] ;
 wire \core.CPU_rd_a2[4] ;
 wire \core.CPU_rd_a3[0] ;
 wire \core.CPU_rd_a3[1] ;
 wire \core.CPU_rd_a3[3] ;
 wire \core.CPU_rd_a3[4] ;
 wire \core.CPU_rd_a4[0] ;
 wire \core.CPU_rd_a4[1] ;
 wire \core.CPU_rd_a4[3] ;
 wire \core.CPU_rd_a4[4] ;
 wire \core.CPU_rd_a5[0] ;
 wire \core.CPU_rd_a5[1] ;
 wire \core.CPU_rd_a5[3] ;
 wire \core.CPU_rd_a5[4] ;
 wire \core.CPU_rd_valid_a1 ;
 wire \core.CPU_rd_valid_a2 ;
 wire \core.CPU_rd_valid_a3 ;
 wire \core.CPU_reset_a1 ;
 wire \core.CPU_reset_a2 ;
 wire \core.CPU_reset_a3 ;
 wire \core.CPU_reset_a4 ;
 wire \core.CPU_result_a3[2] ;
 wire \core.CPU_result_a3[3] ;
 wire \core.CPU_result_a3[4] ;
 wire \core.CPU_result_a3[5] ;
 wire \core.CPU_rf_rd_index1_a2[0] ;
 wire \core.CPU_rf_rd_index1_a2[1] ;
 wire \core.CPU_rf_rd_index1_a2[4] ;
 wire \core.CPU_rf_rd_index2_a2[0] ;
 wire \core.CPU_rf_rd_index2_a2[1] ;
 wire \core.CPU_rf_rd_index2_a2[3] ;
 wire \core.CPU_src1_value_a2[0] ;
 wire \core.CPU_src1_value_a2[10] ;
 wire \core.CPU_src1_value_a2[11] ;
 wire \core.CPU_src1_value_a2[12] ;
 wire \core.CPU_src1_value_a2[13] ;
 wire \core.CPU_src1_value_a2[14] ;
 wire \core.CPU_src1_value_a2[15] ;
 wire \core.CPU_src1_value_a2[16] ;
 wire \core.CPU_src1_value_a2[17] ;
 wire \core.CPU_src1_value_a2[18] ;
 wire \core.CPU_src1_value_a2[19] ;
 wire \core.CPU_src1_value_a2[1] ;
 wire \core.CPU_src1_value_a2[20] ;
 wire \core.CPU_src1_value_a2[21] ;
 wire \core.CPU_src1_value_a2[22] ;
 wire \core.CPU_src1_value_a2[23] ;
 wire \core.CPU_src1_value_a2[24] ;
 wire \core.CPU_src1_value_a2[25] ;
 wire \core.CPU_src1_value_a2[26] ;
 wire \core.CPU_src1_value_a2[27] ;
 wire \core.CPU_src1_value_a2[28] ;
 wire \core.CPU_src1_value_a2[29] ;
 wire \core.CPU_src1_value_a2[2] ;
 wire \core.CPU_src1_value_a2[30] ;
 wire \core.CPU_src1_value_a2[31] ;
 wire \core.CPU_src1_value_a2[3] ;
 wire \core.CPU_src1_value_a2[4] ;
 wire \core.CPU_src1_value_a2[5] ;
 wire \core.CPU_src1_value_a2[6] ;
 wire \core.CPU_src1_value_a2[7] ;
 wire \core.CPU_src1_value_a2[8] ;
 wire \core.CPU_src1_value_a2[9] ;
 wire \core.CPU_src1_value_a3[0] ;
 wire \core.CPU_src1_value_a3[10] ;
 wire \core.CPU_src1_value_a3[11] ;
 wire \core.CPU_src1_value_a3[12] ;
 wire \core.CPU_src1_value_a3[13] ;
 wire \core.CPU_src1_value_a3[14] ;
 wire \core.CPU_src1_value_a3[15] ;
 wire \core.CPU_src1_value_a3[16] ;
 wire \core.CPU_src1_value_a3[17] ;
 wire \core.CPU_src1_value_a3[18] ;
 wire \core.CPU_src1_value_a3[19] ;
 wire \core.CPU_src1_value_a3[1] ;
 wire \core.CPU_src1_value_a3[20] ;
 wire \core.CPU_src1_value_a3[21] ;
 wire \core.CPU_src1_value_a3[22] ;
 wire \core.CPU_src1_value_a3[23] ;
 wire \core.CPU_src1_value_a3[24] ;
 wire \core.CPU_src1_value_a3[25] ;
 wire \core.CPU_src1_value_a3[26] ;
 wire \core.CPU_src1_value_a3[27] ;
 wire \core.CPU_src1_value_a3[28] ;
 wire \core.CPU_src1_value_a3[29] ;
 wire \core.CPU_src1_value_a3[2] ;
 wire \core.CPU_src1_value_a3[30] ;
 wire \core.CPU_src1_value_a3[31] ;
 wire \core.CPU_src1_value_a3[3] ;
 wire \core.CPU_src1_value_a3[4] ;
 wire \core.CPU_src1_value_a3[5] ;
 wire \core.CPU_src1_value_a3[6] ;
 wire \core.CPU_src1_value_a3[7] ;
 wire \core.CPU_src1_value_a3[8] ;
 wire \core.CPU_src1_value_a3[9] ;
 wire \core.CPU_src2_value_a2[0] ;
 wire \core.CPU_src2_value_a2[10] ;
 wire \core.CPU_src2_value_a2[11] ;
 wire \core.CPU_src2_value_a2[12] ;
 wire \core.CPU_src2_value_a2[13] ;
 wire \core.CPU_src2_value_a2[14] ;
 wire \core.CPU_src2_value_a2[15] ;
 wire \core.CPU_src2_value_a2[16] ;
 wire \core.CPU_src2_value_a2[17] ;
 wire \core.CPU_src2_value_a2[18] ;
 wire \core.CPU_src2_value_a2[19] ;
 wire \core.CPU_src2_value_a2[1] ;
 wire \core.CPU_src2_value_a2[20] ;
 wire \core.CPU_src2_value_a2[21] ;
 wire \core.CPU_src2_value_a2[22] ;
 wire \core.CPU_src2_value_a2[23] ;
 wire \core.CPU_src2_value_a2[24] ;
 wire \core.CPU_src2_value_a2[25] ;
 wire \core.CPU_src2_value_a2[26] ;
 wire \core.CPU_src2_value_a2[27] ;
 wire \core.CPU_src2_value_a2[28] ;
 wire \core.CPU_src2_value_a2[29] ;
 wire \core.CPU_src2_value_a2[2] ;
 wire \core.CPU_src2_value_a2[30] ;
 wire \core.CPU_src2_value_a2[31] ;
 wire \core.CPU_src2_value_a2[3] ;
 wire \core.CPU_src2_value_a2[4] ;
 wire \core.CPU_src2_value_a2[5] ;
 wire \core.CPU_src2_value_a2[6] ;
 wire \core.CPU_src2_value_a2[7] ;
 wire \core.CPU_src2_value_a2[8] ;
 wire \core.CPU_src2_value_a2[9] ;
 wire \core.CPU_src2_value_a3[0] ;
 wire \core.CPU_src2_value_a3[10] ;
 wire \core.CPU_src2_value_a3[11] ;
 wire \core.CPU_src2_value_a3[12] ;
 wire \core.CPU_src2_value_a3[13] ;
 wire \core.CPU_src2_value_a3[14] ;
 wire \core.CPU_src2_value_a3[15] ;
 wire \core.CPU_src2_value_a3[16] ;
 wire \core.CPU_src2_value_a3[17] ;
 wire \core.CPU_src2_value_a3[18] ;
 wire \core.CPU_src2_value_a3[19] ;
 wire \core.CPU_src2_value_a3[1] ;
 wire \core.CPU_src2_value_a3[20] ;
 wire \core.CPU_src2_value_a3[21] ;
 wire \core.CPU_src2_value_a3[22] ;
 wire \core.CPU_src2_value_a3[23] ;
 wire \core.CPU_src2_value_a3[24] ;
 wire \core.CPU_src2_value_a3[25] ;
 wire \core.CPU_src2_value_a3[26] ;
 wire \core.CPU_src2_value_a3[27] ;
 wire \core.CPU_src2_value_a3[28] ;
 wire \core.CPU_src2_value_a3[29] ;
 wire \core.CPU_src2_value_a3[2] ;
 wire \core.CPU_src2_value_a3[30] ;
 wire \core.CPU_src2_value_a3[31] ;
 wire \core.CPU_src2_value_a3[3] ;
 wire \core.CPU_src2_value_a3[4] ;
 wire \core.CPU_src2_value_a3[5] ;
 wire \core.CPU_src2_value_a3[6] ;
 wire \core.CPU_src2_value_a3[7] ;
 wire \core.CPU_src2_value_a3[8] ;
 wire \core.CPU_src2_value_a3[9] ;
 wire \core.CPU_valid_a4 ;
 wire \core.CPU_valid_load_a3 ;
 wire \core.CPU_valid_load_a5 ;
 wire \core.CPU_valid_taken_br_a4 ;
 wire \core.CPU_valid_taken_br_a5 ;
 wire \core.w_CPU_dmem_rd_data_a4[0] ;
 wire \core.w_CPU_dmem_rd_data_a4[10] ;
 wire \core.w_CPU_dmem_rd_data_a4[11] ;
 wire \core.w_CPU_dmem_rd_data_a4[12] ;
 wire \core.w_CPU_dmem_rd_data_a4[13] ;
 wire \core.w_CPU_dmem_rd_data_a4[14] ;
 wire \core.w_CPU_dmem_rd_data_a4[15] ;
 wire \core.w_CPU_dmem_rd_data_a4[16] ;
 wire \core.w_CPU_dmem_rd_data_a4[17] ;
 wire \core.w_CPU_dmem_rd_data_a4[18] ;
 wire \core.w_CPU_dmem_rd_data_a4[19] ;
 wire \core.w_CPU_dmem_rd_data_a4[1] ;
 wire \core.w_CPU_dmem_rd_data_a4[20] ;
 wire \core.w_CPU_dmem_rd_data_a4[21] ;
 wire \core.w_CPU_dmem_rd_data_a4[22] ;
 wire \core.w_CPU_dmem_rd_data_a4[23] ;
 wire \core.w_CPU_dmem_rd_data_a4[24] ;
 wire \core.w_CPU_dmem_rd_data_a4[25] ;
 wire \core.w_CPU_dmem_rd_data_a4[26] ;
 wire \core.w_CPU_dmem_rd_data_a4[27] ;
 wire \core.w_CPU_dmem_rd_data_a4[28] ;
 wire \core.w_CPU_dmem_rd_data_a4[29] ;
 wire \core.w_CPU_dmem_rd_data_a4[2] ;
 wire \core.w_CPU_dmem_rd_data_a4[30] ;
 wire \core.w_CPU_dmem_rd_data_a4[31] ;
 wire \core.w_CPU_dmem_rd_data_a4[3] ;
 wire \core.w_CPU_dmem_rd_data_a4[4] ;
 wire \core.w_CPU_dmem_rd_data_a4[5] ;
 wire \core.w_CPU_dmem_rd_data_a4[6] ;
 wire \core.w_CPU_dmem_rd_data_a4[7] ;
 wire \core.w_CPU_dmem_rd_data_a4[8] ;
 wire \core.w_CPU_dmem_rd_data_a4[9] ;
 wire net;
 wire net1;
 wire net2;
 wire net3;

 sky130_fd_sc_hd__or4_2 _05430_ (.A(\core.CPU_valid_load_a5 ),
    .B(\core.CPU_valid_taken_br_a5 ),
    .C(\core.CPU_valid_taken_br_a4 ),
    .D(\core.CPU_dmem_rd_en_a4 ),
    .X(_01114_));
 sky130_fd_sc_hd__inv_2 _05431_ (.A(_01114_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2b_1 _05439_ (.A(\core.CPU_is_beq_a3 ),
    .B_N(\core.CPU_is_bne_a3 ),
    .Y(_01122_));
 sky130_fd_sc_hd__nand4_1 _05444_ (.A(_00110_),
    .B(_00116_),
    .C(_00124_),
    .D(_00130_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand2_1 _05447_ (.A(_00136_),
    .B(_00142_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _05450_ (.A(_00148_),
    .B(_00154_),
    .Y(_01133_));
 sky130_fd_sc_hd__nand2_1 _05453_ (.A(_00160_),
    .B(_00166_),
    .Y(_01136_));
 sky130_fd_sc_hd__nor4_1 _05454_ (.A(_01127_),
    .B(_01130_),
    .C(_01133_),
    .D(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__nand4_1 _05459_ (.A(_00086_),
    .B(_00092_),
    .C(_00098_),
    .D(_00104_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand3_1 _05463_ (.A(_00070_),
    .B(_00076_),
    .C(_00080_),
    .Y(_01146_));
 sky130_fd_sc_hd__nand4_1 _05468_ (.A(_00046_),
    .B(_00052_),
    .C(_00056_),
    .D(_00062_),
    .Y(_01151_));
 sky130_fd_sc_hd__nand3_1 _05470_ (.A(_00040_),
    .B(_00034_),
    .C(_00022_),
    .Y(_01153_));
 sky130_fd_sc_hd__nor4_1 _05471_ (.A(_01142_),
    .B(_01146_),
    .C(_01151_),
    .D(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__xor2_1 _05472_ (.A(net585),
    .B(\core.CPU_src1_value_a3[31] ),
    .X(_01155_));
 sky130_fd_sc_hd__and3_1 _05474_ (.A(_00172_),
    .B(_00178_),
    .C(_00184_),
    .X(_01157_));
 sky130_fd_sc_hd__nand2_1 _05476_ (.A(_00029_),
    .B(_01157_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand3_1 _05480_ (.A(_00025_),
    .B(_00194_),
    .C(_00200_),
    .Y(_01163_));
 sky130_fd_sc_hd__nor3_1 _05481_ (.A(_01155_),
    .B(_01159_),
    .C(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__nand3_1 _05482_ (.A(_01137_),
    .B(_01154_),
    .C(_01164_),
    .Y(_01165_));
 sky130_fd_sc_hd__mux2i_1 _05483_ (.A0(\core.CPU_is_beq_a3 ),
    .A1(_01122_),
    .S(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__nor2_1 _05484_ (.A(net562),
    .B(_01166_),
    .Y(_01167_));
 sky130_fd_sc_hd__nand2_1 _05486_ (.A(\core.CPU_is_load_a3 ),
    .B(net536),
    .Y(_01168_));
 sky130_fd_sc_hd__inv_1 _05487_ (.A(_01168_),
    .Y(\core.CPU_valid_load_a3 ));
 sky130_fd_sc_hd__inv_1 _05488_ (.A(\core.CPU_src1_value_a3[0] ),
    .Y(_00021_));
 sky130_fd_sc_hd__inv_1 _05489_ (.A(\core.CPU_src1_value_a3[1] ),
    .Y(_00003_));
 sky130_fd_sc_hd__inv_1 _05490_ (.A(\core.CPU_imem_rd_addr_a1[0] ),
    .Y(\core.CPU_inc_pc_a1[2] ));
 sky130_fd_sc_hd__xor2_1 _05492_ (.A(\core.CPU_imem_rd_addr_a1[2] ),
    .B(_00207_),
    .X(\core.CPU_inc_pc_a1[4] ));
 sky130_fd_sc_hd__nand3_1 _05493_ (.A(\core.CPU_imem_rd_addr_a1[2] ),
    .B(\core.CPU_imem_rd_addr_a1[1] ),
    .C(\core.CPU_imem_rd_addr_a1[0] ),
    .Y(_01170_));
 sky130_fd_sc_hd__xnor2_1 _05494_ (.A(net614),
    .B(_01170_),
    .Y(\core.CPU_inc_pc_a1[5] ));
 sky130_fd_sc_hd__inv_1 _05500_ (.A(_00204_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand2b_1 _05503_ (.A_N(\core.CPU_imem_rd_addr_a1[3] ),
    .B(_00206_),
    .Y(_01179_));
 sky130_fd_sc_hd__nor4_1 _05504_ (.A(net615),
    .B(_00205_),
    .C(_00207_),
    .D(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__a31oi_1 _05505_ (.A1(net615),
    .A2(\core.CPU_imem_rd_addr_a1[3] ),
    .A3(_01176_),
    .B1(_01180_),
    .Y(\core.CPU_imem_rd_data_a1[7] ));
 sky130_fd_sc_hd__nand2b_1 _05506_ (.A_N(\core.CPU_imem_rd_addr_a1[3] ),
    .B(_00205_),
    .Y(_01181_));
 sky130_fd_sc_hd__nor2b_1 _05507_ (.A(_00206_),
    .B_N(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__o21ai_0 _05508_ (.A1(net615),
    .A2(_01182_),
    .B1(_01179_),
    .Y(\core.CPU_imem_rd_data_a1[8] ));
 sky130_fd_sc_hd__nor2_1 _05509_ (.A(_00205_),
    .B(_00206_),
    .Y(_01183_));
 sky130_fd_sc_hd__a21o_1 _05510_ (.A1(_00204_),
    .A2(_01183_),
    .B1(\core.CPU_imem_rd_addr_a1[3] ),
    .X(_01184_));
 sky130_fd_sc_hd__a21oi_1 _05511_ (.A1(\core.CPU_imem_rd_addr_a1[3] ),
    .A2(_00204_),
    .B1(_00207_),
    .Y(_01185_));
 sky130_fd_sc_hd__nor3_1 _05512_ (.A(_00205_),
    .B(_00206_),
    .C(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__a21oi_1 _05513_ (.A1(net615),
    .A2(_01184_),
    .B1(_01186_),
    .Y(\core.CPU_imem_rd_data_a1[10] ));
 sky130_fd_sc_hd__o22a_1 _05514_ (.A1(net615),
    .A2(net614),
    .B1(_00205_),
    .B2(_00204_),
    .X(_01187_));
 sky130_fd_sc_hd__nor2_1 _05515_ (.A(_00207_),
    .B(_01187_),
    .Y(_01188_));
 sky130_fd_sc_hd__a21oi_1 _05516_ (.A1(\core.CPU_imem_rd_addr_a1[2] ),
    .A2(net614),
    .B1(_01188_),
    .Y(\core.CPU_imem_rd_data_a1[11] ));
 sky130_fd_sc_hd__inv_1 _05517_ (.A(\core.CPU_imm_a2[1] ),
    .Y(_00010_));
 sky130_fd_sc_hd__inv_1 _05518_ (.A(\core.CPU_inc_pc_a2[1] ),
    .Y(_00011_));
 sky130_fd_sc_hd__inv_1 _05519_ (.A(_00202_),
    .Y(_00012_));
 sky130_fd_sc_hd__inv_1 _05520_ (.A(_00014_),
    .Y(\core.CPU_br_tgt_pc_a2[1] ));
 sky130_fd_sc_hd__inv_1 _05521_ (.A(\core.CPU_src2_value_a3[28] ),
    .Y(_00023_));
 sky130_fd_sc_hd__inv_1 _05522_ (.A(\core.CPU_src2_value_a3[27] ),
    .Y(_00027_));
 sky130_fd_sc_hd__inv_1 _05523_ (.A(\core.CPU_src2_value_a3[1] ),
    .Y(_00035_));
 sky130_fd_sc_hd__inv_1 _05524_ (.A(\core.CPU_src2_value_a3[2] ),
    .Y(_00038_));
 sky130_fd_sc_hd__inv_1 _05525_ (.A(\core.CPU_src2_value_a3[3] ),
    .Y(_00044_));
 sky130_fd_sc_hd__inv_1 _05526_ (.A(\core.CPU_src2_value_a3[4] ),
    .Y(_00050_));
 sky130_fd_sc_hd__inv_1 _05527_ (.A(\core.CPU_src2_value_a3[5] ),
    .Y(_00054_));
 sky130_fd_sc_hd__inv_1 _05528_ (.A(\core.CPU_src2_value_a3[6] ),
    .Y(_00060_));
 sky130_fd_sc_hd__inv_1 _05529_ (.A(\core.CPU_src2_value_a3[7] ),
    .Y(_00068_));
 sky130_fd_sc_hd__inv_1 _05530_ (.A(\core.CPU_src2_value_a3[8] ),
    .Y(_00074_));
 sky130_fd_sc_hd__inv_1 _05531_ (.A(\core.CPU_src2_value_a3[9] ),
    .Y(_00078_));
 sky130_fd_sc_hd__inv_1 _05532_ (.A(\core.CPU_src2_value_a3[10] ),
    .Y(_00084_));
 sky130_fd_sc_hd__inv_1 _05533_ (.A(\core.CPU_src2_value_a3[11] ),
    .Y(_00090_));
 sky130_fd_sc_hd__inv_1 _05534_ (.A(\core.CPU_src2_value_a3[12] ),
    .Y(_00096_));
 sky130_fd_sc_hd__inv_1 _05535_ (.A(\core.CPU_src2_value_a3[13] ),
    .Y(_00102_));
 sky130_fd_sc_hd__inv_1 _05536_ (.A(\core.CPU_src2_value_a3[14] ),
    .Y(_00108_));
 sky130_fd_sc_hd__inv_1 _05537_ (.A(\core.CPU_src2_value_a3[15] ),
    .Y(_00114_));
 sky130_fd_sc_hd__inv_1 _05538_ (.A(\core.CPU_src2_value_a3[16] ),
    .Y(_00122_));
 sky130_fd_sc_hd__inv_1 _05539_ (.A(\core.CPU_src2_value_a3[17] ),
    .Y(_00128_));
 sky130_fd_sc_hd__inv_1 _05540_ (.A(\core.CPU_src2_value_a3[18] ),
    .Y(_00134_));
 sky130_fd_sc_hd__inv_1 _05541_ (.A(\core.CPU_src2_value_a3[19] ),
    .Y(_00140_));
 sky130_fd_sc_hd__inv_1 _05542_ (.A(\core.CPU_src2_value_a3[20] ),
    .Y(_00146_));
 sky130_fd_sc_hd__inv_1 _05543_ (.A(\core.CPU_src2_value_a3[21] ),
    .Y(_00152_));
 sky130_fd_sc_hd__inv_1 _05544_ (.A(\core.CPU_src2_value_a3[22] ),
    .Y(_00158_));
 sky130_fd_sc_hd__inv_1 _05545_ (.A(\core.CPU_src2_value_a3[23] ),
    .Y(_00164_));
 sky130_fd_sc_hd__inv_1 _05546_ (.A(\core.CPU_src2_value_a3[24] ),
    .Y(_00170_));
 sky130_fd_sc_hd__inv_1 _05547_ (.A(\core.CPU_src2_value_a3[25] ),
    .Y(_00176_));
 sky130_fd_sc_hd__inv_1 _05548_ (.A(\core.CPU_src2_value_a3[26] ),
    .Y(_00182_));
 sky130_fd_sc_hd__inv_1 _05549_ (.A(net586),
    .Y(_00192_));
 sky130_fd_sc_hd__inv_1 _05550_ (.A(\core.CPU_src2_value_a3[30] ),
    .Y(_00198_));
 sky130_fd_sc_hd__inv_1 _05551_ (.A(\core.CPU_imem_rd_addr_a1[1] ),
    .Y(_00203_));
 sky130_fd_sc_hd__nand2_1 _05554_ (.A(\core.CPU_is_s_instr_a4 ),
    .B(\core.CPU_valid_a4 ),
    .Y(_01191_));
 sky130_fd_sc_hd__nor2_1 _05558_ (.A(\core.CPU_dmem_addr_a4[3] ),
    .B(\core.CPU_dmem_addr_a4[2] ),
    .Y(_01195_));
 sky130_fd_sc_hd__nor2_1 _05561_ (.A(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_2 _05562_ (.A(_01195_),
    .B(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hd__nor2_4 _05563_ (.A(net561),
    .B(net534),
    .Y(_01200_));
 sky130_fd_sc_hd__nand2_1 _05565_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(_01200_),
    .Y(_01202_));
 sky130_fd_sc_hd__and2_0 _05566_ (.A(\core.CPU_is_s_instr_a4 ),
    .B(\core.CPU_valid_a4 ),
    .X(_01203_));
 sky130_fd_sc_hd__nor4_2 _05569_ (.A(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .C(\core.CPU_dmem_addr_a4[3] ),
    .D(\core.CPU_dmem_addr_a4[2] ),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_2 _05570_ (.A(net560),
    .B(net558),
    .Y(_01207_));
 sky130_fd_sc_hd__nand2_1 _05572_ (.A(\core.CPU_Dmem_value_a5[0][0] ),
    .B(_01207_),
    .Y(_01209_));
 sky130_fd_sc_hd__a21oi_1 _05576_ (.A1(_01202_),
    .A2(_01209_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _05579_ (.A(net584),
    .B(net457),
    .Y(_01215_));
 sky130_fd_sc_hd__nand2_1 _05580_ (.A(\core.CPU_Dmem_value_a5[0][10] ),
    .B(net533),
    .Y(_01216_));
 sky130_fd_sc_hd__a21oi_1 _05581_ (.A1(_01215_),
    .A2(_01216_),
    .B1(net601),
    .Y(_00209_));
 sky130_fd_sc_hd__nand2_1 _05584_ (.A(net583),
    .B(net457),
    .Y(_01219_));
 sky130_fd_sc_hd__nand2_1 _05585_ (.A(\core.CPU_Dmem_value_a5[0][11] ),
    .B(net533),
    .Y(_01220_));
 sky130_fd_sc_hd__a21oi_1 _05586_ (.A1(_01219_),
    .A2(_01220_),
    .B1(net600),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _05589_ (.A(net582),
    .B(net457),
    .Y(_01223_));
 sky130_fd_sc_hd__nand2_1 _05590_ (.A(\core.CPU_Dmem_value_a5[0][12] ),
    .B(net533),
    .Y(_01224_));
 sky130_fd_sc_hd__a21oi_1 _05591_ (.A1(_01223_),
    .A2(_01224_),
    .B1(net600),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _05594_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net457),
    .Y(_01227_));
 sky130_fd_sc_hd__nand2_1 _05595_ (.A(\core.CPU_Dmem_value_a5[0][13] ),
    .B(net533),
    .Y(_01228_));
 sky130_fd_sc_hd__a21oi_1 _05596_ (.A1(_01227_),
    .A2(_01228_),
    .B1(net604),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _05599_ (.A(net581),
    .B(net457),
    .Y(_01231_));
 sky130_fd_sc_hd__nand2_1 _05600_ (.A(\core.CPU_Dmem_value_a5[0][14] ),
    .B(_01207_),
    .Y(_01232_));
 sky130_fd_sc_hd__a21oi_1 _05601_ (.A1(_01231_),
    .A2(_01232_),
    .B1(net599),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _05604_ (.A(net580),
    .B(net457),
    .Y(_01235_));
 sky130_fd_sc_hd__nand2_1 _05605_ (.A(\core.CPU_Dmem_value_a5[0][15] ),
    .B(net533),
    .Y(_01236_));
 sky130_fd_sc_hd__a21oi_1 _05606_ (.A1(_01235_),
    .A2(_01236_),
    .B1(net603),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _05609_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(_01200_),
    .Y(_01239_));
 sky130_fd_sc_hd__nand2_1 _05610_ (.A(\core.CPU_Dmem_value_a5[0][16] ),
    .B(_01207_),
    .Y(_01240_));
 sky130_fd_sc_hd__a21oi_1 _05611_ (.A1(_01239_),
    .A2(_01240_),
    .B1(net604),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _05614_ (.A(net579),
    .B(net457),
    .Y(_01243_));
 sky130_fd_sc_hd__nand2_1 _05615_ (.A(\core.CPU_Dmem_value_a5[0][17] ),
    .B(net533),
    .Y(_01244_));
 sky130_fd_sc_hd__a21oi_1 _05616_ (.A1(_01243_),
    .A2(_01244_),
    .B1(net604),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _05619_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net457),
    .Y(_01247_));
 sky130_fd_sc_hd__nand2_1 _05620_ (.A(\core.CPU_Dmem_value_a5[0][18] ),
    .B(_01207_),
    .Y(_01248_));
 sky130_fd_sc_hd__a21oi_1 _05621_ (.A1(_01247_),
    .A2(_01248_),
    .B1(net604),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_1 _05625_ (.A(net578),
    .B(net457),
    .Y(_01252_));
 sky130_fd_sc_hd__nand2_1 _05627_ (.A(\core.CPU_Dmem_value_a5[0][19] ),
    .B(_01207_),
    .Y(_01254_));
 sky130_fd_sc_hd__a21oi_1 _05629_ (.A1(_01252_),
    .A2(_01254_),
    .B1(net600),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _05632_ (.A(net577),
    .B(net457),
    .Y(_01258_));
 sky130_fd_sc_hd__nand2_1 _05633_ (.A(\core.CPU_Dmem_value_a5[0][1] ),
    .B(net533),
    .Y(_01259_));
 sky130_fd_sc_hd__a21oi_1 _05634_ (.A1(_01258_),
    .A2(_01259_),
    .B1(net605),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_1 _05637_ (.A(net576),
    .B(net457),
    .Y(_01262_));
 sky130_fd_sc_hd__nand2_1 _05638_ (.A(\core.CPU_Dmem_value_a5[0][20] ),
    .B(_01207_),
    .Y(_01263_));
 sky130_fd_sc_hd__a21oi_1 _05639_ (.A1(_01262_),
    .A2(_01263_),
    .B1(net601),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_1 _05642_ (.A(net575),
    .B(net457),
    .Y(_01266_));
 sky130_fd_sc_hd__nand2_1 _05643_ (.A(\core.CPU_Dmem_value_a5[0][21] ),
    .B(net533),
    .Y(_01267_));
 sky130_fd_sc_hd__a21oi_1 _05644_ (.A1(_01266_),
    .A2(_01267_),
    .B1(net603),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _05647_ (.A(net574),
    .B(net457),
    .Y(_01270_));
 sky130_fd_sc_hd__nand2_1 _05648_ (.A(\core.CPU_Dmem_value_a5[0][22] ),
    .B(net533),
    .Y(_01271_));
 sky130_fd_sc_hd__a21oi_1 _05649_ (.A1(_01270_),
    .A2(_01271_),
    .B1(net601),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_1 _05652_ (.A(net573),
    .B(net457),
    .Y(_01274_));
 sky130_fd_sc_hd__nand2_1 _05653_ (.A(\core.CPU_Dmem_value_a5[0][23] ),
    .B(net533),
    .Y(_01275_));
 sky130_fd_sc_hd__a21oi_1 _05654_ (.A1(_01274_),
    .A2(_01275_),
    .B1(net601),
    .Y(_00223_));
 sky130_fd_sc_hd__nand2_1 _05657_ (.A(net572),
    .B(net457),
    .Y(_01278_));
 sky130_fd_sc_hd__nand2_1 _05658_ (.A(\core.CPU_Dmem_value_a5[0][24] ),
    .B(_01207_),
    .Y(_01279_));
 sky130_fd_sc_hd__a21oi_1 _05659_ (.A1(_01278_),
    .A2(_01279_),
    .B1(net601),
    .Y(_00224_));
 sky130_fd_sc_hd__nand2_1 _05662_ (.A(net571),
    .B(net457),
    .Y(_01282_));
 sky130_fd_sc_hd__nand2_1 _05663_ (.A(\core.CPU_Dmem_value_a5[0][25] ),
    .B(_01207_),
    .Y(_01283_));
 sky130_fd_sc_hd__a21oi_1 _05664_ (.A1(_01282_),
    .A2(_01283_),
    .B1(net600),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_1 _05667_ (.A(net570),
    .B(net457),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _05668_ (.A(\core.CPU_Dmem_value_a5[0][26] ),
    .B(net533),
    .Y(_01287_));
 sky130_fd_sc_hd__a21oi_1 _05669_ (.A1(_01286_),
    .A2(_01287_),
    .B1(net603),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _05672_ (.A(net569),
    .B(net457),
    .Y(_01290_));
 sky130_fd_sc_hd__nand2_1 _05673_ (.A(\core.CPU_Dmem_value_a5[0][27] ),
    .B(net533),
    .Y(_01291_));
 sky130_fd_sc_hd__a21oi_1 _05674_ (.A1(_01290_),
    .A2(_01291_),
    .B1(net604),
    .Y(_00227_));
 sky130_fd_sc_hd__nand2_1 _05678_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net457),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _05680_ (.A(\core.CPU_Dmem_value_a5[0][28] ),
    .B(_01207_),
    .Y(_01297_));
 sky130_fd_sc_hd__a21oi_1 _05682_ (.A1(_01295_),
    .A2(_01297_),
    .B1(net603),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _05685_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net457),
    .Y(_01301_));
 sky130_fd_sc_hd__nand2_1 _05686_ (.A(\core.CPU_Dmem_value_a5[0][29] ),
    .B(net533),
    .Y(_01302_));
 sky130_fd_sc_hd__a21oi_1 _05687_ (.A1(_01301_),
    .A2(_01302_),
    .B1(net599),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _05690_ (.A(net568),
    .B(net457),
    .Y(_01305_));
 sky130_fd_sc_hd__nand2_1 _05691_ (.A(\core.CPU_Dmem_value_a5[0][2] ),
    .B(net533),
    .Y(_01306_));
 sky130_fd_sc_hd__a21oi_1 _05692_ (.A1(_01305_),
    .A2(_01306_),
    .B1(net605),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _05695_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net457),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _05696_ (.A(\core.CPU_Dmem_value_a5[0][30] ),
    .B(_01207_),
    .Y(_01310_));
 sky130_fd_sc_hd__a21oi_1 _05697_ (.A1(_01309_),
    .A2(_01310_),
    .B1(net602),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _05700_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net457),
    .Y(_01313_));
 sky130_fd_sc_hd__nand2_1 _05701_ (.A(\core.CPU_Dmem_value_a5[0][31] ),
    .B(net533),
    .Y(_01314_));
 sky130_fd_sc_hd__a21oi_1 _05702_ (.A1(_01313_),
    .A2(_01314_),
    .B1(net601),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _05705_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net457),
    .Y(_01317_));
 sky130_fd_sc_hd__nand2_1 _05706_ (.A(\core.CPU_Dmem_value_a5[0][3] ),
    .B(_01207_),
    .Y(_01318_));
 sky130_fd_sc_hd__a21oi_1 _05707_ (.A1(_01317_),
    .A2(_01318_),
    .B1(net602),
    .Y(_00233_));
 sky130_fd_sc_hd__nand2_1 _05710_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(_01200_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand2_1 _05711_ (.A(\core.CPU_Dmem_value_a5[0][4] ),
    .B(_01207_),
    .Y(_01322_));
 sky130_fd_sc_hd__a21oi_1 _05712_ (.A1(_01321_),
    .A2(_01322_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _05715_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net457),
    .Y(_01325_));
 sky130_fd_sc_hd__nand2_1 _05716_ (.A(\core.CPU_Dmem_value_a5[0][5] ),
    .B(_01207_),
    .Y(_01326_));
 sky130_fd_sc_hd__a21oi_1 _05717_ (.A1(_01325_),
    .A2(_01326_),
    .B1(net605),
    .Y(_00235_));
 sky130_fd_sc_hd__nand2_1 _05720_ (.A(net567),
    .B(net457),
    .Y(_01329_));
 sky130_fd_sc_hd__nand2_1 _05721_ (.A(\core.CPU_Dmem_value_a5[0][6] ),
    .B(net533),
    .Y(_01330_));
 sky130_fd_sc_hd__a21oi_1 _05722_ (.A1(_01329_),
    .A2(_01330_),
    .B1(net602),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _05725_ (.A(net566),
    .B(net457),
    .Y(_01333_));
 sky130_fd_sc_hd__nand2_1 _05726_ (.A(\core.CPU_Dmem_value_a5[0][7] ),
    .B(net533),
    .Y(_01334_));
 sky130_fd_sc_hd__a21oi_1 _05727_ (.A1(_01333_),
    .A2(_01334_),
    .B1(net602),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _05730_ (.A(net565),
    .B(net457),
    .Y(_01337_));
 sky130_fd_sc_hd__nand2_1 _05731_ (.A(\core.CPU_Dmem_value_a5[0][8] ),
    .B(net533),
    .Y(_01338_));
 sky130_fd_sc_hd__a21oi_1 _05733_ (.A1(_01337_),
    .A2(_01338_),
    .B1(net601),
    .Y(_00238_));
 sky130_fd_sc_hd__nand2_1 _05736_ (.A(net564),
    .B(net457),
    .Y(_01342_));
 sky130_fd_sc_hd__nand2_1 _05737_ (.A(\core.CPU_Dmem_value_a5[0][9] ),
    .B(net533),
    .Y(_01343_));
 sky130_fd_sc_hd__a21oi_1 _05738_ (.A1(_01342_),
    .A2(_01343_),
    .B1(net603),
    .Y(_00239_));
 sky130_fd_sc_hd__nand2b_1 _05739_ (.A_N(\core.CPU_dmem_addr_a4[0] ),
    .B(\core.CPU_dmem_addr_a4[1] ),
    .Y(_01344_));
 sky130_fd_sc_hd__nand2b_1 _05741_ (.A_N(\core.CPU_dmem_addr_a4[2] ),
    .B(\core.CPU_dmem_addr_a4[3] ),
    .Y(_01346_));
 sky130_fd_sc_hd__nor3_2 _05743_ (.A(net561),
    .B(_01344_),
    .C(_01346_),
    .Y(_01348_));
 sky130_fd_sc_hd__nand2_1 _05745_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net532),
    .Y(_01350_));
 sky130_fd_sc_hd__nor2_4 _05746_ (.A(_01344_),
    .B(_01346_),
    .Y(_01351_));
 sky130_fd_sc_hd__nand2_2 _05747_ (.A(net560),
    .B(net529),
    .Y(_01352_));
 sky130_fd_sc_hd__nand2_1 _05749_ (.A(\core.CPU_Dmem_value_a5[10][0] ),
    .B(_01352_),
    .Y(_01354_));
 sky130_fd_sc_hd__a21oi_1 _05750_ (.A1(_01350_),
    .A2(_01354_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _05751_ (.A(net584),
    .B(net531),
    .Y(_01355_));
 sky130_fd_sc_hd__nand2_1 _05752_ (.A(\core.CPU_Dmem_value_a5[10][10] ),
    .B(net456),
    .Y(_01356_));
 sky130_fd_sc_hd__a21oi_1 _05753_ (.A1(_01355_),
    .A2(_01356_),
    .B1(net601),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _05754_ (.A(net583),
    .B(net531),
    .Y(_01357_));
 sky130_fd_sc_hd__nand2_1 _05755_ (.A(\core.CPU_Dmem_value_a5[10][11] ),
    .B(net456),
    .Y(_01358_));
 sky130_fd_sc_hd__a21oi_1 _05756_ (.A1(_01357_),
    .A2(_01358_),
    .B1(net600),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _05757_ (.A(net582),
    .B(net531),
    .Y(_01359_));
 sky130_fd_sc_hd__nand2_1 _05758_ (.A(\core.CPU_Dmem_value_a5[10][12] ),
    .B(net456),
    .Y(_01360_));
 sky130_fd_sc_hd__a21oi_1 _05759_ (.A1(_01359_),
    .A2(_01360_),
    .B1(net602),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _05760_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net532),
    .Y(_01361_));
 sky130_fd_sc_hd__nand2_1 _05761_ (.A(\core.CPU_Dmem_value_a5[10][13] ),
    .B(net456),
    .Y(_01362_));
 sky130_fd_sc_hd__a21oi_1 _05762_ (.A1(_01361_),
    .A2(_01362_),
    .B1(net605),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _05763_ (.A(net581),
    .B(net531),
    .Y(_01363_));
 sky130_fd_sc_hd__nand2_1 _05764_ (.A(\core.CPU_Dmem_value_a5[10][14] ),
    .B(_01352_),
    .Y(_01364_));
 sky130_fd_sc_hd__a21oi_1 _05765_ (.A1(_01363_),
    .A2(_01364_),
    .B1(net602),
    .Y(_00245_));
 sky130_fd_sc_hd__nand2_1 _05766_ (.A(net580),
    .B(net532),
    .Y(_01365_));
 sky130_fd_sc_hd__nand2_1 _05767_ (.A(\core.CPU_Dmem_value_a5[10][15] ),
    .B(net456),
    .Y(_01366_));
 sky130_fd_sc_hd__a21oi_1 _05768_ (.A1(_01365_),
    .A2(_01366_),
    .B1(net603),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _05769_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net532),
    .Y(_01367_));
 sky130_fd_sc_hd__nand2_1 _05770_ (.A(\core.CPU_Dmem_value_a5[10][16] ),
    .B(_01352_),
    .Y(_01368_));
 sky130_fd_sc_hd__a21oi_1 _05771_ (.A1(_01367_),
    .A2(_01368_),
    .B1(net604),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _05773_ (.A(net579),
    .B(net532),
    .Y(_01370_));
 sky130_fd_sc_hd__nand2_1 _05775_ (.A(\core.CPU_Dmem_value_a5[10][17] ),
    .B(_01352_),
    .Y(_01372_));
 sky130_fd_sc_hd__a21oi_1 _05777_ (.A1(_01370_),
    .A2(_01372_),
    .B1(net604),
    .Y(_00248_));
 sky130_fd_sc_hd__nand2_1 _05778_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net532),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _05779_ (.A(\core.CPU_Dmem_value_a5[10][18] ),
    .B(_01352_),
    .Y(_01375_));
 sky130_fd_sc_hd__a21oi_1 _05780_ (.A1(_01374_),
    .A2(_01375_),
    .B1(net604),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_1 _05781_ (.A(net578),
    .B(net532),
    .Y(_01376_));
 sky130_fd_sc_hd__nand2_1 _05782_ (.A(\core.CPU_Dmem_value_a5[10][19] ),
    .B(net456),
    .Y(_01377_));
 sky130_fd_sc_hd__a21oi_1 _05783_ (.A1(_01376_),
    .A2(_01377_),
    .B1(net600),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _05785_ (.A(\core.CPU_Dmem_value_a5[10][1] ),
    .B(net456),
    .Y(_01379_));
 sky130_fd_sc_hd__nand2_1 _05786_ (.A(net577),
    .B(net532),
    .Y(_01380_));
 sky130_fd_sc_hd__nand3b_1 _05787_ (.A_N(net605),
    .B(_01379_),
    .C(_01380_),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_1 _05788_ (.A(net576),
    .B(net532),
    .Y(_01381_));
 sky130_fd_sc_hd__nand2_1 _05789_ (.A(\core.CPU_Dmem_value_a5[10][20] ),
    .B(net456),
    .Y(_01382_));
 sky130_fd_sc_hd__a21oi_1 _05790_ (.A1(_01381_),
    .A2(_01382_),
    .B1(net601),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _05791_ (.A(net575),
    .B(net532),
    .Y(_01383_));
 sky130_fd_sc_hd__nand2_1 _05792_ (.A(\core.CPU_Dmem_value_a5[10][21] ),
    .B(net456),
    .Y(_01384_));
 sky130_fd_sc_hd__a21oi_1 _05793_ (.A1(_01383_),
    .A2(_01384_),
    .B1(net601),
    .Y(_00253_));
 sky130_fd_sc_hd__nand2_1 _05794_ (.A(net574),
    .B(net531),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_1 _05795_ (.A(\core.CPU_Dmem_value_a5[10][22] ),
    .B(net456),
    .Y(_01386_));
 sky130_fd_sc_hd__a21oi_1 _05796_ (.A1(_01385_),
    .A2(_01386_),
    .B1(net601),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _05797_ (.A(net573),
    .B(net532),
    .Y(_01387_));
 sky130_fd_sc_hd__nand2_1 _05798_ (.A(\core.CPU_Dmem_value_a5[10][23] ),
    .B(net456),
    .Y(_01388_));
 sky130_fd_sc_hd__a21oi_1 _05799_ (.A1(_01387_),
    .A2(_01388_),
    .B1(net601),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _05800_ (.A(net572),
    .B(net532),
    .Y(_01389_));
 sky130_fd_sc_hd__nand2_1 _05801_ (.A(\core.CPU_Dmem_value_a5[10][24] ),
    .B(net456),
    .Y(_01390_));
 sky130_fd_sc_hd__a21oi_1 _05802_ (.A1(_01389_),
    .A2(_01390_),
    .B1(net601),
    .Y(_00256_));
 sky130_fd_sc_hd__nand2_1 _05803_ (.A(net571),
    .B(net532),
    .Y(_01391_));
 sky130_fd_sc_hd__nand2_1 _05804_ (.A(\core.CPU_Dmem_value_a5[10][25] ),
    .B(_01352_),
    .Y(_01392_));
 sky130_fd_sc_hd__a21oi_1 _05805_ (.A1(_01391_),
    .A2(_01392_),
    .B1(net600),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_1 _05806_ (.A(net570),
    .B(net532),
    .Y(_01393_));
 sky130_fd_sc_hd__nand2_1 _05807_ (.A(\core.CPU_Dmem_value_a5[10][26] ),
    .B(net456),
    .Y(_01394_));
 sky130_fd_sc_hd__a21oi_1 _05808_ (.A1(_01393_),
    .A2(_01394_),
    .B1(net603),
    .Y(_00258_));
 sky130_fd_sc_hd__nand2_1 _05810_ (.A(net569),
    .B(net532),
    .Y(_01396_));
 sky130_fd_sc_hd__nand2_1 _05812_ (.A(\core.CPU_Dmem_value_a5[10][27] ),
    .B(_01352_),
    .Y(_01398_));
 sky130_fd_sc_hd__a21oi_1 _05814_ (.A1(_01396_),
    .A2(_01398_),
    .B1(net604),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _05815_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net532),
    .Y(_01400_));
 sky130_fd_sc_hd__nand2_1 _05816_ (.A(\core.CPU_Dmem_value_a5[10][28] ),
    .B(_01352_),
    .Y(_01401_));
 sky130_fd_sc_hd__a21oi_1 _05817_ (.A1(_01400_),
    .A2(_01401_),
    .B1(net603),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _05818_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net531),
    .Y(_01402_));
 sky130_fd_sc_hd__nand2_1 _05819_ (.A(\core.CPU_Dmem_value_a5[10][29] ),
    .B(_01352_),
    .Y(_01403_));
 sky130_fd_sc_hd__a21oi_1 _05820_ (.A1(_01402_),
    .A2(_01403_),
    .B1(net599),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_1 _05821_ (.A(net568),
    .B(net532),
    .Y(_01404_));
 sky130_fd_sc_hd__nand2_1 _05822_ (.A(\core.CPU_Dmem_value_a5[10][2] ),
    .B(net456),
    .Y(_01405_));
 sky130_fd_sc_hd__a21oi_1 _05823_ (.A1(_01404_),
    .A2(_01405_),
    .B1(net605),
    .Y(_00262_));
 sky130_fd_sc_hd__nand2_1 _05824_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net531),
    .Y(_01406_));
 sky130_fd_sc_hd__nand2_1 _05825_ (.A(\core.CPU_Dmem_value_a5[10][30] ),
    .B(_01352_),
    .Y(_01407_));
 sky130_fd_sc_hd__a21oi_1 _05826_ (.A1(_01406_),
    .A2(_01407_),
    .B1(net602),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _05827_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net531),
    .Y(_01408_));
 sky130_fd_sc_hd__nand2_1 _05828_ (.A(\core.CPU_Dmem_value_a5[10][31] ),
    .B(net456),
    .Y(_01409_));
 sky130_fd_sc_hd__a21oi_1 _05829_ (.A1(_01408_),
    .A2(_01409_),
    .B1(net601),
    .Y(_00264_));
 sky130_fd_sc_hd__nand2_1 _05830_ (.A(\core.CPU_Dmem_value_a5[10][3] ),
    .B(_01352_),
    .Y(_01410_));
 sky130_fd_sc_hd__nand2_1 _05831_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net531),
    .Y(_01411_));
 sky130_fd_sc_hd__nand3b_1 _05832_ (.A_N(net599),
    .B(_01410_),
    .C(_01411_),
    .Y(_00265_));
 sky130_fd_sc_hd__nand2_1 _05833_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net532),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _05834_ (.A(\core.CPU_Dmem_value_a5[10][4] ),
    .B(_01352_),
    .Y(_01413_));
 sky130_fd_sc_hd__a21oi_1 _05835_ (.A1(_01412_),
    .A2(_01413_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00266_));
 sky130_fd_sc_hd__nand2_1 _05836_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net532),
    .Y(_01414_));
 sky130_fd_sc_hd__nand2_1 _05837_ (.A(\core.CPU_Dmem_value_a5[10][5] ),
    .B(net456),
    .Y(_01415_));
 sky130_fd_sc_hd__a21oi_1 _05838_ (.A1(_01414_),
    .A2(_01415_),
    .B1(net605),
    .Y(_00267_));
 sky130_fd_sc_hd__nand2_1 _05839_ (.A(net567),
    .B(net531),
    .Y(_01416_));
 sky130_fd_sc_hd__nand2_1 _05840_ (.A(\core.CPU_Dmem_value_a5[10][6] ),
    .B(net456),
    .Y(_01417_));
 sky130_fd_sc_hd__a21oi_1 _05841_ (.A1(_01416_),
    .A2(_01417_),
    .B1(net599),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _05842_ (.A(net566),
    .B(net531),
    .Y(_01418_));
 sky130_fd_sc_hd__nand2_1 _05843_ (.A(\core.CPU_Dmem_value_a5[10][7] ),
    .B(net456),
    .Y(_01419_));
 sky130_fd_sc_hd__a21oi_1 _05844_ (.A1(_01418_),
    .A2(_01419_),
    .B1(net602),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _05845_ (.A(net565),
    .B(net531),
    .Y(_01420_));
 sky130_fd_sc_hd__nand2_1 _05846_ (.A(\core.CPU_Dmem_value_a5[10][8] ),
    .B(net456),
    .Y(_01421_));
 sky130_fd_sc_hd__a21oi_1 _05848_ (.A1(_01420_),
    .A2(_01421_),
    .B1(net601),
    .Y(_00270_));
 sky130_fd_sc_hd__nand2_1 _05849_ (.A(net564),
    .B(net532),
    .Y(_01423_));
 sky130_fd_sc_hd__nand2_1 _05850_ (.A(\core.CPU_Dmem_value_a5[10][9] ),
    .B(net456),
    .Y(_01424_));
 sky130_fd_sc_hd__a21oi_1 _05851_ (.A1(_01423_),
    .A2(_01424_),
    .B1(net603),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _05852_ (.A(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .Y(_01425_));
 sky130_fd_sc_hd__nor2_4 _05853_ (.A(_01346_),
    .B(_01425_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_2 _05854_ (.A(net560),
    .B(net527),
    .Y(_01427_));
 sky130_fd_sc_hd__nand2_1 _05856_ (.A(\core.CPU_Dmem_value_a5[11][0] ),
    .B(_01427_),
    .Y(_01429_));
 sky130_fd_sc_hd__nor3_2 _05857_ (.A(net561),
    .B(_01346_),
    .C(_01425_),
    .Y(_01430_));
 sky130_fd_sc_hd__nand2_1 _05859_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net526),
    .Y(_01432_));
 sky130_fd_sc_hd__nand3b_1 _05860_ (.A_N(\core.CPU_reset_a4 ),
    .B(_01429_),
    .C(_01432_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand2_1 _05861_ (.A(net584),
    .B(net526),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _05862_ (.A(\core.CPU_Dmem_value_a5[11][10] ),
    .B(net455),
    .Y(_01434_));
 sky130_fd_sc_hd__a21oi_1 _05863_ (.A1(_01433_),
    .A2(_01434_),
    .B1(net601),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _05864_ (.A(net583),
    .B(net526),
    .Y(_01435_));
 sky130_fd_sc_hd__nand2_1 _05865_ (.A(\core.CPU_Dmem_value_a5[11][11] ),
    .B(net455),
    .Y(_01436_));
 sky130_fd_sc_hd__a21oi_1 _05866_ (.A1(_01435_),
    .A2(_01436_),
    .B1(net600),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _05867_ (.A(net582),
    .B(net526),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_1 _05868_ (.A(\core.CPU_Dmem_value_a5[11][12] ),
    .B(net455),
    .Y(_01438_));
 sky130_fd_sc_hd__a21oi_1 _05869_ (.A1(_01437_),
    .A2(_01438_),
    .B1(net600),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2_1 _05870_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net526),
    .Y(_01439_));
 sky130_fd_sc_hd__nand2_1 _05871_ (.A(\core.CPU_Dmem_value_a5[11][13] ),
    .B(net455),
    .Y(_01440_));
 sky130_fd_sc_hd__a21oi_1 _05872_ (.A1(_01439_),
    .A2(_01440_),
    .B1(net605),
    .Y(_00276_));
 sky130_fd_sc_hd__nand2_1 _05873_ (.A(net581),
    .B(net526),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_1 _05874_ (.A(\core.CPU_Dmem_value_a5[11][14] ),
    .B(_01427_),
    .Y(_01442_));
 sky130_fd_sc_hd__a21oi_1 _05875_ (.A1(_01441_),
    .A2(_01442_),
    .B1(net602),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _05876_ (.A(net580),
    .B(net526),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_1 _05877_ (.A(\core.CPU_Dmem_value_a5[11][15] ),
    .B(net455),
    .Y(_01444_));
 sky130_fd_sc_hd__a21oi_1 _05878_ (.A1(_01443_),
    .A2(_01444_),
    .B1(net603),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _05879_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net526),
    .Y(_01445_));
 sky130_fd_sc_hd__nand2_1 _05880_ (.A(\core.CPU_Dmem_value_a5[11][16] ),
    .B(_01427_),
    .Y(_01446_));
 sky130_fd_sc_hd__a21oi_1 _05881_ (.A1(_01445_),
    .A2(_01446_),
    .B1(net603),
    .Y(_00279_));
 sky130_fd_sc_hd__nand2_1 _05883_ (.A(net579),
    .B(net526),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_1 _05885_ (.A(\core.CPU_Dmem_value_a5[11][17] ),
    .B(net455),
    .Y(_01450_));
 sky130_fd_sc_hd__a21oi_1 _05886_ (.A1(_01448_),
    .A2(_01450_),
    .B1(net604),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _05887_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net526),
    .Y(_01451_));
 sky130_fd_sc_hd__nand2_1 _05888_ (.A(\core.CPU_Dmem_value_a5[11][18] ),
    .B(_01427_),
    .Y(_01452_));
 sky130_fd_sc_hd__a21oi_1 _05890_ (.A1(_01451_),
    .A2(_01452_),
    .B1(net604),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_1 _05891_ (.A(net578),
    .B(net526),
    .Y(_01454_));
 sky130_fd_sc_hd__nand2_1 _05892_ (.A(\core.CPU_Dmem_value_a5[11][19] ),
    .B(_01427_),
    .Y(_01455_));
 sky130_fd_sc_hd__a21oi_1 _05893_ (.A1(_01454_),
    .A2(_01455_),
    .B1(net600),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2_1 _05894_ (.A(\core.CPU_Dmem_value_a5[11][1] ),
    .B(net455),
    .Y(_01456_));
 sky130_fd_sc_hd__nand2_1 _05895_ (.A(net577),
    .B(net526),
    .Y(_01457_));
 sky130_fd_sc_hd__nand3b_1 _05896_ (.A_N(net605),
    .B(_01456_),
    .C(_01457_),
    .Y(_00283_));
 sky130_fd_sc_hd__nand2_1 _05897_ (.A(net576),
    .B(net526),
    .Y(_01458_));
 sky130_fd_sc_hd__nand2_1 _05898_ (.A(\core.CPU_Dmem_value_a5[11][20] ),
    .B(_01427_),
    .Y(_01459_));
 sky130_fd_sc_hd__a21oi_1 _05899_ (.A1(_01458_),
    .A2(_01459_),
    .B1(net601),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _05900_ (.A(net575),
    .B(net526),
    .Y(_01460_));
 sky130_fd_sc_hd__nand2_1 _05901_ (.A(\core.CPU_Dmem_value_a5[11][21] ),
    .B(net455),
    .Y(_01461_));
 sky130_fd_sc_hd__a21oi_1 _05902_ (.A1(_01460_),
    .A2(_01461_),
    .B1(net605),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _05903_ (.A(net574),
    .B(net526),
    .Y(_01462_));
 sky130_fd_sc_hd__nand2_1 _05904_ (.A(\core.CPU_Dmem_value_a5[11][22] ),
    .B(net455),
    .Y(_01463_));
 sky130_fd_sc_hd__a21oi_1 _05905_ (.A1(_01462_),
    .A2(_01463_),
    .B1(net601),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_1 _05906_ (.A(net573),
    .B(net526),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2_1 _05907_ (.A(\core.CPU_Dmem_value_a5[11][23] ),
    .B(net455),
    .Y(_01465_));
 sky130_fd_sc_hd__a21oi_1 _05908_ (.A1(_01464_),
    .A2(_01465_),
    .B1(net601),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_1 _05909_ (.A(net572),
    .B(net526),
    .Y(_01466_));
 sky130_fd_sc_hd__nand2_1 _05910_ (.A(\core.CPU_Dmem_value_a5[11][24] ),
    .B(net455),
    .Y(_01467_));
 sky130_fd_sc_hd__a21oi_1 _05911_ (.A1(_01466_),
    .A2(_01467_),
    .B1(net600),
    .Y(_00288_));
 sky130_fd_sc_hd__nand2_1 _05912_ (.A(net571),
    .B(net526),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _05913_ (.A(\core.CPU_Dmem_value_a5[11][25] ),
    .B(_01427_),
    .Y(_01469_));
 sky130_fd_sc_hd__a21oi_1 _05914_ (.A1(_01468_),
    .A2(_01469_),
    .B1(net600),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _05915_ (.A(net570),
    .B(net526),
    .Y(_01470_));
 sky130_fd_sc_hd__nand2_1 _05916_ (.A(\core.CPU_Dmem_value_a5[11][26] ),
    .B(_01427_),
    .Y(_01471_));
 sky130_fd_sc_hd__a21oi_1 _05917_ (.A1(_01470_),
    .A2(_01471_),
    .B1(net603),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _05919_ (.A(net569),
    .B(net526),
    .Y(_01473_));
 sky130_fd_sc_hd__nand2_1 _05921_ (.A(\core.CPU_Dmem_value_a5[11][27] ),
    .B(net455),
    .Y(_01475_));
 sky130_fd_sc_hd__a21oi_1 _05922_ (.A1(_01473_),
    .A2(_01475_),
    .B1(net604),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_1 _05923_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net526),
    .Y(_01476_));
 sky130_fd_sc_hd__nand2_1 _05924_ (.A(\core.CPU_Dmem_value_a5[11][28] ),
    .B(_01427_),
    .Y(_01477_));
 sky130_fd_sc_hd__a21oi_1 _05927_ (.A1(_01476_),
    .A2(_01477_),
    .B1(net600),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _05928_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net526),
    .Y(_01480_));
 sky130_fd_sc_hd__nand2_1 _05929_ (.A(\core.CPU_Dmem_value_a5[11][29] ),
    .B(_01427_),
    .Y(_01481_));
 sky130_fd_sc_hd__a21oi_1 _05930_ (.A1(_01480_),
    .A2(_01481_),
    .B1(net602),
    .Y(_00293_));
 sky130_fd_sc_hd__nand2_1 _05931_ (.A(net568),
    .B(net526),
    .Y(_01482_));
 sky130_fd_sc_hd__nand2_1 _05932_ (.A(\core.CPU_Dmem_value_a5[11][2] ),
    .B(net455),
    .Y(_01483_));
 sky130_fd_sc_hd__a21oi_1 _05933_ (.A1(_01482_),
    .A2(_01483_),
    .B1(net605),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _05934_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net526),
    .Y(_01484_));
 sky130_fd_sc_hd__nand2_1 _05935_ (.A(\core.CPU_Dmem_value_a5[11][30] ),
    .B(_01427_),
    .Y(_01485_));
 sky130_fd_sc_hd__a21oi_1 _05936_ (.A1(_01484_),
    .A2(_01485_),
    .B1(net602),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _05937_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net526),
    .Y(_01486_));
 sky130_fd_sc_hd__nand2_1 _05938_ (.A(\core.CPU_Dmem_value_a5[11][31] ),
    .B(net455),
    .Y(_01487_));
 sky130_fd_sc_hd__a21oi_1 _05939_ (.A1(_01486_),
    .A2(_01487_),
    .B1(net601),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _05940_ (.A(\core.CPU_Dmem_value_a5[11][3] ),
    .B(_01427_),
    .Y(_01488_));
 sky130_fd_sc_hd__nand2_1 _05941_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net526),
    .Y(_01489_));
 sky130_fd_sc_hd__nand3b_1 _05942_ (.A_N(net600),
    .B(_01488_),
    .C(_01489_),
    .Y(_00297_));
 sky130_fd_sc_hd__nand2_1 _05943_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net526),
    .Y(_01490_));
 sky130_fd_sc_hd__nand2_1 _05944_ (.A(\core.CPU_Dmem_value_a5[11][4] ),
    .B(_01427_),
    .Y(_01491_));
 sky130_fd_sc_hd__a21oi_1 _05945_ (.A1(_01490_),
    .A2(_01491_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00298_));
 sky130_fd_sc_hd__nand2_1 _05946_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net526),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_1 _05947_ (.A(\core.CPU_Dmem_value_a5[11][5] ),
    .B(_01427_),
    .Y(_01493_));
 sky130_fd_sc_hd__a21oi_1 _05948_ (.A1(_01492_),
    .A2(_01493_),
    .B1(net605),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _05949_ (.A(net567),
    .B(net526),
    .Y(_01494_));
 sky130_fd_sc_hd__nand2_1 _05950_ (.A(\core.CPU_Dmem_value_a5[11][6] ),
    .B(net455),
    .Y(_01495_));
 sky130_fd_sc_hd__a21oi_1 _05951_ (.A1(_01494_),
    .A2(_01495_),
    .B1(net602),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _05952_ (.A(net566),
    .B(net526),
    .Y(_01496_));
 sky130_fd_sc_hd__nand2_1 _05953_ (.A(\core.CPU_Dmem_value_a5[11][7] ),
    .B(net455),
    .Y(_01497_));
 sky130_fd_sc_hd__a21oi_1 _05954_ (.A1(_01496_),
    .A2(_01497_),
    .B1(net602),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _05955_ (.A(net565),
    .B(net526),
    .Y(_01498_));
 sky130_fd_sc_hd__nand2_1 _05956_ (.A(\core.CPU_Dmem_value_a5[11][8] ),
    .B(net455),
    .Y(_01499_));
 sky130_fd_sc_hd__a21oi_1 _05957_ (.A1(_01498_),
    .A2(_01499_),
    .B1(net601),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _05958_ (.A(net564),
    .B(net526),
    .Y(_01500_));
 sky130_fd_sc_hd__nand2_1 _05959_ (.A(\core.CPU_Dmem_value_a5[11][9] ),
    .B(net455),
    .Y(_01501_));
 sky130_fd_sc_hd__a21oi_1 _05961_ (.A1(_01500_),
    .A2(_01501_),
    .B1(net605),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _05962_ (.A(\core.CPU_dmem_addr_a4[3] ),
    .B(\core.CPU_dmem_addr_a4[2] ),
    .Y(_01503_));
 sky130_fd_sc_hd__nor4_2 _05963_ (.A(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .C(net561),
    .D(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__nand2_1 _05965_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net525),
    .Y(_01506_));
 sky130_fd_sc_hd__nor3_2 _05966_ (.A(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .C(_01503_),
    .Y(_01507_));
 sky130_fd_sc_hd__nand2_2 _05967_ (.A(net560),
    .B(net523),
    .Y(_01508_));
 sky130_fd_sc_hd__nand2_1 _05969_ (.A(\core.CPU_Dmem_value_a5[12][0] ),
    .B(net454),
    .Y(_01510_));
 sky130_fd_sc_hd__a21oi_1 _05970_ (.A1(_01506_),
    .A2(_01510_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _05971_ (.A(net584),
    .B(net525),
    .Y(_01511_));
 sky130_fd_sc_hd__nand2_1 _05972_ (.A(\core.CPU_Dmem_value_a5[12][10] ),
    .B(net454),
    .Y(_01512_));
 sky130_fd_sc_hd__a21oi_1 _05973_ (.A1(_01511_),
    .A2(_01512_),
    .B1(net601),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _05974_ (.A(net583),
    .B(net525),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_1 _05975_ (.A(\core.CPU_Dmem_value_a5[12][11] ),
    .B(net454),
    .Y(_01514_));
 sky130_fd_sc_hd__a21oi_1 _05976_ (.A1(_01513_),
    .A2(_01514_),
    .B1(net600),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _05977_ (.A(net582),
    .B(net525),
    .Y(_01515_));
 sky130_fd_sc_hd__nand2_1 _05978_ (.A(\core.CPU_Dmem_value_a5[12][12] ),
    .B(net454),
    .Y(_01516_));
 sky130_fd_sc_hd__a21oi_1 _05979_ (.A1(_01515_),
    .A2(_01516_),
    .B1(net602),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_1 _05980_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net525),
    .Y(_01517_));
 sky130_fd_sc_hd__nand2_1 _05981_ (.A(\core.CPU_Dmem_value_a5[12][13] ),
    .B(net454),
    .Y(_01518_));
 sky130_fd_sc_hd__a21oi_1 _05982_ (.A1(_01517_),
    .A2(_01518_),
    .B1(net604),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _05983_ (.A(net581),
    .B(net525),
    .Y(_01519_));
 sky130_fd_sc_hd__nand2_1 _05984_ (.A(\core.CPU_Dmem_value_a5[12][14] ),
    .B(net454),
    .Y(_01520_));
 sky130_fd_sc_hd__a21oi_1 _05985_ (.A1(_01519_),
    .A2(_01520_),
    .B1(net602),
    .Y(_00309_));
 sky130_fd_sc_hd__nand2_1 _05986_ (.A(net580),
    .B(net525),
    .Y(_01521_));
 sky130_fd_sc_hd__nand2_1 _05987_ (.A(\core.CPU_Dmem_value_a5[12][15] ),
    .B(net454),
    .Y(_01522_));
 sky130_fd_sc_hd__a21oi_1 _05988_ (.A1(_01521_),
    .A2(_01522_),
    .B1(net601),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _05989_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net525),
    .Y(_01523_));
 sky130_fd_sc_hd__nand2_1 _05990_ (.A(\core.CPU_Dmem_value_a5[12][16] ),
    .B(net454),
    .Y(_01524_));
 sky130_fd_sc_hd__a21oi_1 _05991_ (.A1(_01523_),
    .A2(_01524_),
    .B1(net603),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _05993_ (.A(net579),
    .B(net525),
    .Y(_01526_));
 sky130_fd_sc_hd__nand2_1 _05995_ (.A(\core.CPU_Dmem_value_a5[12][17] ),
    .B(net454),
    .Y(_01528_));
 sky130_fd_sc_hd__a21oi_1 _05996_ (.A1(_01526_),
    .A2(_01528_),
    .B1(net604),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _05997_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net525),
    .Y(_01529_));
 sky130_fd_sc_hd__nand2_1 _05998_ (.A(\core.CPU_Dmem_value_a5[12][18] ),
    .B(net454),
    .Y(_01530_));
 sky130_fd_sc_hd__a21oi_1 _06000_ (.A1(_01529_),
    .A2(_01530_),
    .B1(net604),
    .Y(_00313_));
 sky130_fd_sc_hd__nand2_1 _06001_ (.A(net578),
    .B(net525),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _06002_ (.A(\core.CPU_Dmem_value_a5[12][19] ),
    .B(net454),
    .Y(_01533_));
 sky130_fd_sc_hd__a21oi_1 _06003_ (.A1(_01532_),
    .A2(_01533_),
    .B1(net600),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _06004_ (.A(net577),
    .B(net525),
    .Y(_01534_));
 sky130_fd_sc_hd__nand2_1 _06005_ (.A(\core.CPU_Dmem_value_a5[12][1] ),
    .B(net454),
    .Y(_01535_));
 sky130_fd_sc_hd__a21oi_1 _06006_ (.A1(_01534_),
    .A2(_01535_),
    .B1(net605),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_1 _06007_ (.A(net576),
    .B(net525),
    .Y(_01536_));
 sky130_fd_sc_hd__nand2_1 _06008_ (.A(\core.CPU_Dmem_value_a5[12][20] ),
    .B(net454),
    .Y(_01537_));
 sky130_fd_sc_hd__a21oi_1 _06009_ (.A1(_01536_),
    .A2(_01537_),
    .B1(net601),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _06010_ (.A(net575),
    .B(net525),
    .Y(_01538_));
 sky130_fd_sc_hd__nand2_1 _06011_ (.A(\core.CPU_Dmem_value_a5[12][21] ),
    .B(net454),
    .Y(_01539_));
 sky130_fd_sc_hd__a21oi_1 _06012_ (.A1(_01538_),
    .A2(_01539_),
    .B1(net605),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _06013_ (.A(net574),
    .B(net525),
    .Y(_01540_));
 sky130_fd_sc_hd__nand2_1 _06014_ (.A(\core.CPU_Dmem_value_a5[12][22] ),
    .B(net454),
    .Y(_01541_));
 sky130_fd_sc_hd__a21oi_1 _06015_ (.A1(_01540_),
    .A2(_01541_),
    .B1(net601),
    .Y(_00318_));
 sky130_fd_sc_hd__nand2_1 _06016_ (.A(net573),
    .B(net525),
    .Y(_01542_));
 sky130_fd_sc_hd__nand2_1 _06017_ (.A(\core.CPU_Dmem_value_a5[12][23] ),
    .B(net454),
    .Y(_01543_));
 sky130_fd_sc_hd__a21oi_1 _06018_ (.A1(_01542_),
    .A2(_01543_),
    .B1(net601),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _06019_ (.A(net572),
    .B(net525),
    .Y(_01544_));
 sky130_fd_sc_hd__nand2_1 _06020_ (.A(\core.CPU_Dmem_value_a5[12][24] ),
    .B(net454),
    .Y(_01545_));
 sky130_fd_sc_hd__a21oi_1 _06021_ (.A1(_01544_),
    .A2(_01545_),
    .B1(net601),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _06022_ (.A(net571),
    .B(net525),
    .Y(_01546_));
 sky130_fd_sc_hd__nand2_1 _06023_ (.A(\core.CPU_Dmem_value_a5[12][25] ),
    .B(net454),
    .Y(_01547_));
 sky130_fd_sc_hd__a21oi_1 _06024_ (.A1(_01546_),
    .A2(_01547_),
    .B1(net600),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_1 _06026_ (.A(net570),
    .B(net525),
    .Y(_01549_));
 sky130_fd_sc_hd__nand2_1 _06028_ (.A(\core.CPU_Dmem_value_a5[12][26] ),
    .B(net454),
    .Y(_01551_));
 sky130_fd_sc_hd__a21oi_1 _06029_ (.A1(_01549_),
    .A2(_01551_),
    .B1(net603),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _06030_ (.A(net569),
    .B(net525),
    .Y(_01552_));
 sky130_fd_sc_hd__nand2_1 _06031_ (.A(\core.CPU_Dmem_value_a5[12][27] ),
    .B(net454),
    .Y(_01553_));
 sky130_fd_sc_hd__a21oi_1 _06033_ (.A1(_01552_),
    .A2(_01553_),
    .B1(net604),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _06034_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net525),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_1 _06035_ (.A(\core.CPU_Dmem_value_a5[12][28] ),
    .B(net454),
    .Y(_01556_));
 sky130_fd_sc_hd__a21oi_1 _06036_ (.A1(_01555_),
    .A2(_01556_),
    .B1(net600),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _06037_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net525),
    .Y(_01557_));
 sky130_fd_sc_hd__nand2_1 _06038_ (.A(\core.CPU_Dmem_value_a5[12][29] ),
    .B(net454),
    .Y(_01558_));
 sky130_fd_sc_hd__a21oi_1 _06039_ (.A1(_01557_),
    .A2(_01558_),
    .B1(net602),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _06040_ (.A(\core.CPU_Dmem_value_a5[12][2] ),
    .B(net454),
    .Y(_01559_));
 sky130_fd_sc_hd__nand2_1 _06041_ (.A(net568),
    .B(net525),
    .Y(_01560_));
 sky130_fd_sc_hd__nand3b_1 _06042_ (.A_N(net605),
    .B(_01559_),
    .C(_01560_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _06043_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net525),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_1 _06044_ (.A(\core.CPU_Dmem_value_a5[12][30] ),
    .B(net454),
    .Y(_01562_));
 sky130_fd_sc_hd__a21oi_1 _06045_ (.A1(_01561_),
    .A2(_01562_),
    .B1(net602),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _06046_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net525),
    .Y(_01563_));
 sky130_fd_sc_hd__nand2_1 _06047_ (.A(\core.CPU_Dmem_value_a5[12][31] ),
    .B(net454),
    .Y(_01564_));
 sky130_fd_sc_hd__a21oi_1 _06048_ (.A1(_01563_),
    .A2(_01564_),
    .B1(net601),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _06049_ (.A(\core.CPU_Dmem_value_a5[12][3] ),
    .B(net454),
    .Y(_01565_));
 sky130_fd_sc_hd__nand2_1 _06050_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net525),
    .Y(_01566_));
 sky130_fd_sc_hd__nand3b_1 _06051_ (.A_N(net602),
    .B(_01565_),
    .C(_01566_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _06052_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net525),
    .Y(_01567_));
 sky130_fd_sc_hd__nand2_1 _06053_ (.A(\core.CPU_Dmem_value_a5[12][4] ),
    .B(net454),
    .Y(_01568_));
 sky130_fd_sc_hd__a21oi_1 _06054_ (.A1(_01567_),
    .A2(_01568_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _06055_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net525),
    .Y(_01569_));
 sky130_fd_sc_hd__nand2_1 _06056_ (.A(\core.CPU_Dmem_value_a5[12][5] ),
    .B(net454),
    .Y(_01570_));
 sky130_fd_sc_hd__a21oi_1 _06057_ (.A1(_01569_),
    .A2(_01570_),
    .B1(net605),
    .Y(_00331_));
 sky130_fd_sc_hd__nand2_1 _06058_ (.A(net567),
    .B(net525),
    .Y(_01571_));
 sky130_fd_sc_hd__nand2_1 _06059_ (.A(\core.CPU_Dmem_value_a5[12][6] ),
    .B(net454),
    .Y(_01572_));
 sky130_fd_sc_hd__a21oi_1 _06060_ (.A1(_01571_),
    .A2(_01572_),
    .B1(net602),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _06061_ (.A(net566),
    .B(net525),
    .Y(_01573_));
 sky130_fd_sc_hd__nand2_1 _06062_ (.A(\core.CPU_Dmem_value_a5[12][7] ),
    .B(net454),
    .Y(_01574_));
 sky130_fd_sc_hd__a21oi_1 _06063_ (.A1(_01573_),
    .A2(_01574_),
    .B1(net602),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _06064_ (.A(net565),
    .B(net525),
    .Y(_01575_));
 sky130_fd_sc_hd__nand2_1 _06065_ (.A(\core.CPU_Dmem_value_a5[12][8] ),
    .B(net454),
    .Y(_01576_));
 sky130_fd_sc_hd__a21oi_1 _06066_ (.A1(_01575_),
    .A2(_01576_),
    .B1(net601),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _06067_ (.A(net564),
    .B(net525),
    .Y(_01577_));
 sky130_fd_sc_hd__nand2_1 _06068_ (.A(\core.CPU_Dmem_value_a5[12][9] ),
    .B(net454),
    .Y(_01578_));
 sky130_fd_sc_hd__a21oi_1 _06070_ (.A1(_01577_),
    .A2(_01578_),
    .B1(net603),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2b_1 _06071_ (.A_N(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .Y(_01580_));
 sky130_fd_sc_hd__nor2_4 _06073_ (.A(_01503_),
    .B(_01580_),
    .Y(_01582_));
 sky130_fd_sc_hd__nand2_2 _06074_ (.A(net560),
    .B(net522),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _06076_ (.A(\core.CPU_Dmem_value_a5[13][0] ),
    .B(_01583_),
    .Y(_01585_));
 sky130_fd_sc_hd__nor3_2 _06077_ (.A(net561),
    .B(_01503_),
    .C(_01580_),
    .Y(_01586_));
 sky130_fd_sc_hd__nand2_1 _06079_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net521),
    .Y(_01588_));
 sky130_fd_sc_hd__nand3b_1 _06080_ (.A_N(\core.CPU_reset_a4 ),
    .B(_01585_),
    .C(_01588_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _06081_ (.A(net584),
    .B(net521),
    .Y(_01589_));
 sky130_fd_sc_hd__nand2_1 _06082_ (.A(\core.CPU_Dmem_value_a5[13][10] ),
    .B(net453),
    .Y(_01590_));
 sky130_fd_sc_hd__a21oi_1 _06083_ (.A1(_01589_),
    .A2(_01590_),
    .B1(net601),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _06084_ (.A(net583),
    .B(net521),
    .Y(_01591_));
 sky130_fd_sc_hd__nand2_1 _06085_ (.A(\core.CPU_Dmem_value_a5[13][11] ),
    .B(net453),
    .Y(_01592_));
 sky130_fd_sc_hd__a21oi_1 _06086_ (.A1(_01591_),
    .A2(_01592_),
    .B1(net600),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _06087_ (.A(net582),
    .B(net521),
    .Y(_01593_));
 sky130_fd_sc_hd__nand2_1 _06088_ (.A(\core.CPU_Dmem_value_a5[13][12] ),
    .B(net453),
    .Y(_01594_));
 sky130_fd_sc_hd__a21oi_1 _06089_ (.A1(_01593_),
    .A2(_01594_),
    .B1(net602),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _06090_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net521),
    .Y(_01595_));
 sky130_fd_sc_hd__nand2_1 _06091_ (.A(\core.CPU_Dmem_value_a5[13][13] ),
    .B(net453),
    .Y(_01596_));
 sky130_fd_sc_hd__a21oi_1 _06092_ (.A1(_01595_),
    .A2(_01596_),
    .B1(net605),
    .Y(_00340_));
 sky130_fd_sc_hd__nand2_1 _06093_ (.A(net581),
    .B(net521),
    .Y(_01597_));
 sky130_fd_sc_hd__nand2_1 _06094_ (.A(\core.CPU_Dmem_value_a5[13][14] ),
    .B(_01583_),
    .Y(_01598_));
 sky130_fd_sc_hd__a21oi_1 _06095_ (.A1(_01597_),
    .A2(_01598_),
    .B1(net602),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_1 _06096_ (.A(net580),
    .B(net521),
    .Y(_01599_));
 sky130_fd_sc_hd__nand2_1 _06097_ (.A(\core.CPU_Dmem_value_a5[13][15] ),
    .B(net453),
    .Y(_01600_));
 sky130_fd_sc_hd__a21oi_1 _06098_ (.A1(_01599_),
    .A2(_01600_),
    .B1(net603),
    .Y(_00342_));
 sky130_fd_sc_hd__nand2_1 _06099_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net521),
    .Y(_01601_));
 sky130_fd_sc_hd__nand2_1 _06100_ (.A(\core.CPU_Dmem_value_a5[13][16] ),
    .B(_01583_),
    .Y(_01602_));
 sky130_fd_sc_hd__a21oi_1 _06101_ (.A1(_01601_),
    .A2(_01602_),
    .B1(net603),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _06103_ (.A(net579),
    .B(net521),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_1 _06105_ (.A(\core.CPU_Dmem_value_a5[13][17] ),
    .B(net453),
    .Y(_01606_));
 sky130_fd_sc_hd__a21oi_1 _06106_ (.A1(_01604_),
    .A2(_01606_),
    .B1(net604),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_1 _06107_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net521),
    .Y(_01607_));
 sky130_fd_sc_hd__nand2_1 _06108_ (.A(\core.CPU_Dmem_value_a5[13][18] ),
    .B(net453),
    .Y(_01608_));
 sky130_fd_sc_hd__a21oi_1 _06109_ (.A1(_01607_),
    .A2(_01608_),
    .B1(net604),
    .Y(_00345_));
 sky130_fd_sc_hd__nand2_1 _06110_ (.A(net578),
    .B(net521),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_1 _06111_ (.A(\core.CPU_Dmem_value_a5[13][19] ),
    .B(_01583_),
    .Y(_01610_));
 sky130_fd_sc_hd__a21oi_1 _06113_ (.A1(_01609_),
    .A2(_01610_),
    .B1(net600),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _06114_ (.A(net577),
    .B(net521),
    .Y(_01612_));
 sky130_fd_sc_hd__nand2_1 _06115_ (.A(\core.CPU_Dmem_value_a5[13][1] ),
    .B(net453),
    .Y(_01613_));
 sky130_fd_sc_hd__a21oi_1 _06116_ (.A1(_01612_),
    .A2(_01613_),
    .B1(net605),
    .Y(_00347_));
 sky130_fd_sc_hd__nand2_1 _06117_ (.A(net576),
    .B(net521),
    .Y(_01614_));
 sky130_fd_sc_hd__nand2_1 _06118_ (.A(\core.CPU_Dmem_value_a5[13][20] ),
    .B(net453),
    .Y(_01615_));
 sky130_fd_sc_hd__a21oi_1 _06119_ (.A1(_01614_),
    .A2(_01615_),
    .B1(net601),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _06120_ (.A(net575),
    .B(net521),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_1 _06121_ (.A(\core.CPU_Dmem_value_a5[13][21] ),
    .B(net453),
    .Y(_01617_));
 sky130_fd_sc_hd__a21oi_1 _06122_ (.A1(_01616_),
    .A2(_01617_),
    .B1(net605),
    .Y(_00349_));
 sky130_fd_sc_hd__nand2_1 _06123_ (.A(net574),
    .B(net521),
    .Y(_01618_));
 sky130_fd_sc_hd__nand2_1 _06124_ (.A(\core.CPU_Dmem_value_a5[13][22] ),
    .B(net453),
    .Y(_01619_));
 sky130_fd_sc_hd__a21oi_1 _06125_ (.A1(_01618_),
    .A2(_01619_),
    .B1(net601),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _06126_ (.A(net573),
    .B(net521),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_1 _06127_ (.A(\core.CPU_Dmem_value_a5[13][23] ),
    .B(net453),
    .Y(_01621_));
 sky130_fd_sc_hd__a21oi_1 _06128_ (.A1(_01620_),
    .A2(_01621_),
    .B1(net601),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_1 _06129_ (.A(net572),
    .B(net521),
    .Y(_01622_));
 sky130_fd_sc_hd__nand2_1 _06130_ (.A(\core.CPU_Dmem_value_a5[13][24] ),
    .B(net453),
    .Y(_01623_));
 sky130_fd_sc_hd__a21oi_1 _06131_ (.A1(_01622_),
    .A2(_01623_),
    .B1(net601),
    .Y(_00352_));
 sky130_fd_sc_hd__nand2_1 _06132_ (.A(net571),
    .B(net521),
    .Y(_01624_));
 sky130_fd_sc_hd__nand2_1 _06133_ (.A(\core.CPU_Dmem_value_a5[13][25] ),
    .B(_01583_),
    .Y(_01625_));
 sky130_fd_sc_hd__a21oi_1 _06134_ (.A1(_01624_),
    .A2(_01625_),
    .B1(net600),
    .Y(_00353_));
 sky130_fd_sc_hd__nand2_1 _06136_ (.A(net570),
    .B(net521),
    .Y(_01627_));
 sky130_fd_sc_hd__nand2_1 _06138_ (.A(\core.CPU_Dmem_value_a5[13][26] ),
    .B(net453),
    .Y(_01629_));
 sky130_fd_sc_hd__a21oi_1 _06139_ (.A1(_01627_),
    .A2(_01629_),
    .B1(net603),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_1 _06140_ (.A(net569),
    .B(net521),
    .Y(_01630_));
 sky130_fd_sc_hd__nand2_1 _06141_ (.A(\core.CPU_Dmem_value_a5[13][27] ),
    .B(net453),
    .Y(_01631_));
 sky130_fd_sc_hd__a21oi_1 _06142_ (.A1(_01630_),
    .A2(_01631_),
    .B1(net604),
    .Y(_00355_));
 sky130_fd_sc_hd__nand2_1 _06143_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net521),
    .Y(_01632_));
 sky130_fd_sc_hd__nand2_1 _06144_ (.A(\core.CPU_Dmem_value_a5[13][28] ),
    .B(net453),
    .Y(_01633_));
 sky130_fd_sc_hd__a21oi_1 _06146_ (.A1(_01632_),
    .A2(_01633_),
    .B1(net600),
    .Y(_00356_));
 sky130_fd_sc_hd__nand2_1 _06147_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net521),
    .Y(_01635_));
 sky130_fd_sc_hd__nand2_1 _06148_ (.A(\core.CPU_Dmem_value_a5[13][29] ),
    .B(_01583_),
    .Y(_01636_));
 sky130_fd_sc_hd__a21oi_1 _06149_ (.A1(_01635_),
    .A2(_01636_),
    .B1(net602),
    .Y(_00357_));
 sky130_fd_sc_hd__nand2_1 _06150_ (.A(\core.CPU_Dmem_value_a5[13][2] ),
    .B(net453),
    .Y(_01637_));
 sky130_fd_sc_hd__nand2_1 _06151_ (.A(net568),
    .B(net521),
    .Y(_01638_));
 sky130_fd_sc_hd__nand3b_1 _06152_ (.A_N(net605),
    .B(_01637_),
    .C(_01638_),
    .Y(_00358_));
 sky130_fd_sc_hd__nand2_1 _06153_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net521),
    .Y(_01639_));
 sky130_fd_sc_hd__nand2_1 _06154_ (.A(\core.CPU_Dmem_value_a5[13][30] ),
    .B(_01583_),
    .Y(_01640_));
 sky130_fd_sc_hd__a21oi_1 _06155_ (.A1(_01639_),
    .A2(_01640_),
    .B1(net602),
    .Y(_00359_));
 sky130_fd_sc_hd__nand2_1 _06156_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net521),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_1 _06157_ (.A(\core.CPU_Dmem_value_a5[13][31] ),
    .B(net453),
    .Y(_01642_));
 sky130_fd_sc_hd__a21oi_1 _06158_ (.A1(_01641_),
    .A2(_01642_),
    .B1(net601),
    .Y(_00360_));
 sky130_fd_sc_hd__nand2_1 _06159_ (.A(\core.CPU_Dmem_value_a5[13][3] ),
    .B(_01583_),
    .Y(_01643_));
 sky130_fd_sc_hd__nand2_1 _06160_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net521),
    .Y(_01644_));
 sky130_fd_sc_hd__nand3b_1 _06161_ (.A_N(\core.CPU_reset_a4 ),
    .B(_01643_),
    .C(_01644_),
    .Y(_00361_));
 sky130_fd_sc_hd__nand2_1 _06162_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net521),
    .Y(_01645_));
 sky130_fd_sc_hd__nand2_1 _06163_ (.A(\core.CPU_Dmem_value_a5[13][4] ),
    .B(_01583_),
    .Y(_01646_));
 sky130_fd_sc_hd__a21oi_1 _06164_ (.A1(_01645_),
    .A2(_01646_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_1 _06165_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net521),
    .Y(_01647_));
 sky130_fd_sc_hd__nand2_1 _06166_ (.A(\core.CPU_Dmem_value_a5[13][5] ),
    .B(net453),
    .Y(_01648_));
 sky130_fd_sc_hd__a21oi_1 _06167_ (.A1(_01647_),
    .A2(_01648_),
    .B1(net605),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_1 _06168_ (.A(net567),
    .B(net521),
    .Y(_01649_));
 sky130_fd_sc_hd__nand2_1 _06169_ (.A(\core.CPU_Dmem_value_a5[13][6] ),
    .B(_01583_),
    .Y(_01650_));
 sky130_fd_sc_hd__a21oi_1 _06170_ (.A1(_01649_),
    .A2(_01650_),
    .B1(net602),
    .Y(_00364_));
 sky130_fd_sc_hd__nand2_1 _06171_ (.A(net566),
    .B(net521),
    .Y(_01651_));
 sky130_fd_sc_hd__nand2_1 _06172_ (.A(\core.CPU_Dmem_value_a5[13][7] ),
    .B(_01583_),
    .Y(_01652_));
 sky130_fd_sc_hd__a21oi_1 _06173_ (.A1(_01651_),
    .A2(_01652_),
    .B1(net602),
    .Y(_00365_));
 sky130_fd_sc_hd__nand2_1 _06174_ (.A(net565),
    .B(net521),
    .Y(_01653_));
 sky130_fd_sc_hd__nand2_1 _06175_ (.A(\core.CPU_Dmem_value_a5[13][8] ),
    .B(net453),
    .Y(_01654_));
 sky130_fd_sc_hd__a21oi_1 _06176_ (.A1(_01653_),
    .A2(_01654_),
    .B1(net601),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2_1 _06177_ (.A(net564),
    .B(net521),
    .Y(_01655_));
 sky130_fd_sc_hd__nand2_1 _06178_ (.A(\core.CPU_Dmem_value_a5[13][9] ),
    .B(net453),
    .Y(_01656_));
 sky130_fd_sc_hd__a21oi_1 _06179_ (.A1(_01655_),
    .A2(_01656_),
    .B1(net605),
    .Y(_00367_));
 sky130_fd_sc_hd__nor3_2 _06180_ (.A(net561),
    .B(_01344_),
    .C(_01503_),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _06182_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net519),
    .Y(_01659_));
 sky130_fd_sc_hd__nor2_4 _06183_ (.A(_01344_),
    .B(_01503_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_2 _06184_ (.A(net560),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_1 _06186_ (.A(\core.CPU_Dmem_value_a5[14][0] ),
    .B(_01661_),
    .Y(_01663_));
 sky130_fd_sc_hd__a21oi_1 _06188_ (.A1(_01659_),
    .A2(_01663_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00368_));
 sky130_fd_sc_hd__nand2_1 _06189_ (.A(net584),
    .B(net520),
    .Y(_01665_));
 sky130_fd_sc_hd__nand2_1 _06190_ (.A(\core.CPU_Dmem_value_a5[14][10] ),
    .B(net452),
    .Y(_01666_));
 sky130_fd_sc_hd__a21oi_1 _06191_ (.A1(_01665_),
    .A2(_01666_),
    .B1(net601),
    .Y(_00369_));
 sky130_fd_sc_hd__nand2_1 _06192_ (.A(net583),
    .B(net520),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _06193_ (.A(\core.CPU_Dmem_value_a5[14][11] ),
    .B(net452),
    .Y(_01668_));
 sky130_fd_sc_hd__a21oi_1 _06194_ (.A1(_01667_),
    .A2(_01668_),
    .B1(net600),
    .Y(_00370_));
 sky130_fd_sc_hd__nand2_1 _06195_ (.A(net582),
    .B(net520),
    .Y(_01669_));
 sky130_fd_sc_hd__nand2_1 _06196_ (.A(\core.CPU_Dmem_value_a5[14][12] ),
    .B(_01661_),
    .Y(_01670_));
 sky130_fd_sc_hd__a21oi_1 _06197_ (.A1(_01669_),
    .A2(_01670_),
    .B1(net602),
    .Y(_00371_));
 sky130_fd_sc_hd__nand2_1 _06198_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net519),
    .Y(_01671_));
 sky130_fd_sc_hd__nand2_1 _06199_ (.A(\core.CPU_Dmem_value_a5[14][13] ),
    .B(net452),
    .Y(_01672_));
 sky130_fd_sc_hd__a21oi_1 _06200_ (.A1(_01671_),
    .A2(_01672_),
    .B1(net605),
    .Y(_00372_));
 sky130_fd_sc_hd__nand2_1 _06201_ (.A(net581),
    .B(net520),
    .Y(_01673_));
 sky130_fd_sc_hd__nand2_1 _06202_ (.A(\core.CPU_Dmem_value_a5[14][14] ),
    .B(_01661_),
    .Y(_01674_));
 sky130_fd_sc_hd__a21oi_1 _06203_ (.A1(_01673_),
    .A2(_01674_),
    .B1(net599),
    .Y(_00373_));
 sky130_fd_sc_hd__nand2_1 _06204_ (.A(net580),
    .B(net520),
    .Y(_01675_));
 sky130_fd_sc_hd__nand2_1 _06205_ (.A(\core.CPU_Dmem_value_a5[14][15] ),
    .B(net452),
    .Y(_01676_));
 sky130_fd_sc_hd__a21oi_1 _06206_ (.A1(_01675_),
    .A2(_01676_),
    .B1(net603),
    .Y(_00374_));
 sky130_fd_sc_hd__nand2_1 _06208_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net519),
    .Y(_01678_));
 sky130_fd_sc_hd__nand2_1 _06210_ (.A(\core.CPU_Dmem_value_a5[14][16] ),
    .B(_01661_),
    .Y(_01680_));
 sky130_fd_sc_hd__a21oi_1 _06211_ (.A1(_01678_),
    .A2(_01680_),
    .B1(net603),
    .Y(_00375_));
 sky130_fd_sc_hd__nand2_1 _06212_ (.A(net579),
    .B(net519),
    .Y(_01681_));
 sky130_fd_sc_hd__nand2_1 _06213_ (.A(\core.CPU_Dmem_value_a5[14][17] ),
    .B(net452),
    .Y(_01682_));
 sky130_fd_sc_hd__a21oi_1 _06214_ (.A1(_01681_),
    .A2(_01682_),
    .B1(net604),
    .Y(_00376_));
 sky130_fd_sc_hd__nand2_1 _06215_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net519),
    .Y(_01683_));
 sky130_fd_sc_hd__nand2_1 _06216_ (.A(\core.CPU_Dmem_value_a5[14][18] ),
    .B(net452),
    .Y(_01684_));
 sky130_fd_sc_hd__a21oi_1 _06217_ (.A1(_01683_),
    .A2(_01684_),
    .B1(net604),
    .Y(_00377_));
 sky130_fd_sc_hd__nand2_1 _06218_ (.A(net578),
    .B(net520),
    .Y(_01685_));
 sky130_fd_sc_hd__nand2_1 _06219_ (.A(\core.CPU_Dmem_value_a5[14][19] ),
    .B(_01661_),
    .Y(_01686_));
 sky130_fd_sc_hd__a21oi_1 _06221_ (.A1(_01685_),
    .A2(_01686_),
    .B1(net600),
    .Y(_00378_));
 sky130_fd_sc_hd__nand2_1 _06223_ (.A(\core.CPU_Dmem_value_a5[14][1] ),
    .B(net452),
    .Y(_01689_));
 sky130_fd_sc_hd__nand2_1 _06224_ (.A(net577),
    .B(net519),
    .Y(_01690_));
 sky130_fd_sc_hd__nand3b_1 _06225_ (.A_N(net605),
    .B(_01689_),
    .C(_01690_),
    .Y(_00379_));
 sky130_fd_sc_hd__nand2_1 _06226_ (.A(net576),
    .B(net520),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _06227_ (.A(\core.CPU_Dmem_value_a5[14][20] ),
    .B(_01661_),
    .Y(_01692_));
 sky130_fd_sc_hd__a21oi_1 _06228_ (.A1(_01691_),
    .A2(_01692_),
    .B1(net601),
    .Y(_00380_));
 sky130_fd_sc_hd__nand2_1 _06229_ (.A(net575),
    .B(net520),
    .Y(_01693_));
 sky130_fd_sc_hd__nand2_1 _06230_ (.A(\core.CPU_Dmem_value_a5[14][21] ),
    .B(net452),
    .Y(_01694_));
 sky130_fd_sc_hd__a21oi_1 _06231_ (.A1(_01693_),
    .A2(_01694_),
    .B1(net601),
    .Y(_00381_));
 sky130_fd_sc_hd__nand2_1 _06232_ (.A(net574),
    .B(net520),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _06233_ (.A(\core.CPU_Dmem_value_a5[14][22] ),
    .B(net452),
    .Y(_01696_));
 sky130_fd_sc_hd__a21oi_1 _06234_ (.A1(_01695_),
    .A2(_01696_),
    .B1(net601),
    .Y(_00382_));
 sky130_fd_sc_hd__nand2_1 _06235_ (.A(net573),
    .B(net520),
    .Y(_01697_));
 sky130_fd_sc_hd__nand2_1 _06236_ (.A(\core.CPU_Dmem_value_a5[14][23] ),
    .B(net452),
    .Y(_01698_));
 sky130_fd_sc_hd__a21oi_1 _06237_ (.A1(_01697_),
    .A2(_01698_),
    .B1(net601),
    .Y(_00383_));
 sky130_fd_sc_hd__nand2_1 _06238_ (.A(net572),
    .B(net520),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_1 _06239_ (.A(\core.CPU_Dmem_value_a5[14][24] ),
    .B(_01661_),
    .Y(_01700_));
 sky130_fd_sc_hd__a21oi_1 _06240_ (.A1(_01699_),
    .A2(_01700_),
    .B1(net600),
    .Y(_00384_));
 sky130_fd_sc_hd__nand2_1 _06241_ (.A(net571),
    .B(net520),
    .Y(_01701_));
 sky130_fd_sc_hd__nand2_1 _06242_ (.A(\core.CPU_Dmem_value_a5[14][25] ),
    .B(_01661_),
    .Y(_01702_));
 sky130_fd_sc_hd__a21oi_1 _06243_ (.A1(_01701_),
    .A2(_01702_),
    .B1(net600),
    .Y(_00385_));
 sky130_fd_sc_hd__nand2_1 _06245_ (.A(net570),
    .B(net520),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_1 _06247_ (.A(\core.CPU_Dmem_value_a5[14][26] ),
    .B(net452),
    .Y(_01706_));
 sky130_fd_sc_hd__a21oi_1 _06248_ (.A1(_01704_),
    .A2(_01706_),
    .B1(net603),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _06249_ (.A(net569),
    .B(net519),
    .Y(_01707_));
 sky130_fd_sc_hd__nand2_1 _06250_ (.A(\core.CPU_Dmem_value_a5[14][27] ),
    .B(net452),
    .Y(_01708_));
 sky130_fd_sc_hd__a21oi_1 _06251_ (.A1(_01707_),
    .A2(_01708_),
    .B1(net604),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _06252_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net520),
    .Y(_01709_));
 sky130_fd_sc_hd__nand2_1 _06253_ (.A(\core.CPU_Dmem_value_a5[14][28] ),
    .B(net452),
    .Y(_01710_));
 sky130_fd_sc_hd__a21oi_1 _06254_ (.A1(_01709_),
    .A2(_01710_),
    .B1(net603),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _06255_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net520),
    .Y(_01711_));
 sky130_fd_sc_hd__nand2_1 _06256_ (.A(\core.CPU_Dmem_value_a5[14][29] ),
    .B(_01661_),
    .Y(_01712_));
 sky130_fd_sc_hd__a21oi_1 _06258_ (.A1(_01711_),
    .A2(_01712_),
    .B1(net599),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _06259_ (.A(\core.CPU_Dmem_value_a5[14][2] ),
    .B(net452),
    .Y(_01714_));
 sky130_fd_sc_hd__nand2_1 _06260_ (.A(net568),
    .B(net520),
    .Y(_01715_));
 sky130_fd_sc_hd__nand3b_1 _06261_ (.A_N(net605),
    .B(_01714_),
    .C(_01715_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _06262_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net520),
    .Y(_01716_));
 sky130_fd_sc_hd__nand2_1 _06263_ (.A(\core.CPU_Dmem_value_a5[14][30] ),
    .B(_01661_),
    .Y(_01717_));
 sky130_fd_sc_hd__a21oi_1 _06264_ (.A1(_01716_),
    .A2(_01717_),
    .B1(net599),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_1 _06265_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net520),
    .Y(_01718_));
 sky130_fd_sc_hd__nand2_1 _06266_ (.A(\core.CPU_Dmem_value_a5[14][31] ),
    .B(net452),
    .Y(_01719_));
 sky130_fd_sc_hd__a21oi_1 _06267_ (.A1(_01718_),
    .A2(_01719_),
    .B1(net601),
    .Y(_00392_));
 sky130_fd_sc_hd__nand2_1 _06268_ (.A(\core.CPU_Dmem_value_a5[14][3] ),
    .B(_01661_),
    .Y(_01720_));
 sky130_fd_sc_hd__nand2_1 _06269_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net520),
    .Y(_01721_));
 sky130_fd_sc_hd__nand3b_1 _06270_ (.A_N(net599),
    .B(_01720_),
    .C(_01721_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand2_1 _06271_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net519),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2_1 _06272_ (.A(\core.CPU_Dmem_value_a5[14][4] ),
    .B(_01661_),
    .Y(_01723_));
 sky130_fd_sc_hd__a21oi_1 _06273_ (.A1(_01722_),
    .A2(_01723_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_1 _06274_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net520),
    .Y(_01724_));
 sky130_fd_sc_hd__nand2_1 _06275_ (.A(\core.CPU_Dmem_value_a5[14][5] ),
    .B(net452),
    .Y(_01725_));
 sky130_fd_sc_hd__a21oi_1 _06276_ (.A1(_01724_),
    .A2(_01725_),
    .B1(net605),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _06277_ (.A(net567),
    .B(net520),
    .Y(_01726_));
 sky130_fd_sc_hd__nand2_1 _06278_ (.A(\core.CPU_Dmem_value_a5[14][6] ),
    .B(_01661_),
    .Y(_01727_));
 sky130_fd_sc_hd__a21oi_1 _06279_ (.A1(_01726_),
    .A2(_01727_),
    .B1(net599),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_1 _06280_ (.A(net566),
    .B(net520),
    .Y(_01728_));
 sky130_fd_sc_hd__nand2_1 _06281_ (.A(\core.CPU_Dmem_value_a5[14][7] ),
    .B(_01661_),
    .Y(_01729_));
 sky130_fd_sc_hd__a21oi_1 _06282_ (.A1(_01728_),
    .A2(_01729_),
    .B1(net602),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_1 _06283_ (.A(net565),
    .B(net520),
    .Y(_01730_));
 sky130_fd_sc_hd__nand2_1 _06284_ (.A(\core.CPU_Dmem_value_a5[14][8] ),
    .B(net452),
    .Y(_01731_));
 sky130_fd_sc_hd__a21oi_1 _06285_ (.A1(_01730_),
    .A2(_01731_),
    .B1(net601),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _06286_ (.A(net564),
    .B(net520),
    .Y(_01732_));
 sky130_fd_sc_hd__nand2_1 _06287_ (.A(\core.CPU_Dmem_value_a5[14][9] ),
    .B(net452),
    .Y(_01733_));
 sky130_fd_sc_hd__a21oi_1 _06288_ (.A1(_01732_),
    .A2(_01733_),
    .B1(net605),
    .Y(_00399_));
 sky130_fd_sc_hd__nor2_4 _06289_ (.A(_01425_),
    .B(_01503_),
    .Y(_01734_));
 sky130_fd_sc_hd__nand2_2 _06290_ (.A(net560),
    .B(net517),
    .Y(_01735_));
 sky130_fd_sc_hd__nand2_1 _06292_ (.A(\core.CPU_Dmem_value_a5[15][0] ),
    .B(net451),
    .Y(_01737_));
 sky130_fd_sc_hd__nor3_2 _06293_ (.A(net561),
    .B(_01425_),
    .C(_01503_),
    .Y(_01738_));
 sky130_fd_sc_hd__nand2_1 _06295_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net515),
    .Y(_01740_));
 sky130_fd_sc_hd__nand3b_1 _06296_ (.A_N(\core.CPU_reset_a4 ),
    .B(_01737_),
    .C(_01740_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2_1 _06297_ (.A(net584),
    .B(net516),
    .Y(_01741_));
 sky130_fd_sc_hd__nand2_1 _06298_ (.A(\core.CPU_Dmem_value_a5[15][10] ),
    .B(net451),
    .Y(_01742_));
 sky130_fd_sc_hd__a21oi_1 _06299_ (.A1(_01741_),
    .A2(_01742_),
    .B1(net601),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _06300_ (.A(net583),
    .B(net516),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_1 _06301_ (.A(\core.CPU_Dmem_value_a5[15][11] ),
    .B(_01735_),
    .Y(_01744_));
 sky130_fd_sc_hd__a21oi_1 _06304_ (.A1(_01743_),
    .A2(_01744_),
    .B1(net600),
    .Y(_00402_));
 sky130_fd_sc_hd__nand2_1 _06305_ (.A(net582),
    .B(net516),
    .Y(_01747_));
 sky130_fd_sc_hd__nand2_1 _06306_ (.A(\core.CPU_Dmem_value_a5[15][12] ),
    .B(_01735_),
    .Y(_01748_));
 sky130_fd_sc_hd__a21oi_1 _06307_ (.A1(_01747_),
    .A2(_01748_),
    .B1(net602),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _06308_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net515),
    .Y(_01749_));
 sky130_fd_sc_hd__nand2_1 _06309_ (.A(\core.CPU_Dmem_value_a5[15][13] ),
    .B(net451),
    .Y(_01750_));
 sky130_fd_sc_hd__a21oi_1 _06310_ (.A1(_01749_),
    .A2(_01750_),
    .B1(net605),
    .Y(_00404_));
 sky130_fd_sc_hd__nand2_1 _06311_ (.A(net581),
    .B(net516),
    .Y(_01751_));
 sky130_fd_sc_hd__nand2_1 _06312_ (.A(\core.CPU_Dmem_value_a5[15][14] ),
    .B(_01735_),
    .Y(_01752_));
 sky130_fd_sc_hd__a21oi_1 _06313_ (.A1(_01751_),
    .A2(_01752_),
    .B1(net602),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _06314_ (.A(net580),
    .B(net516),
    .Y(_01753_));
 sky130_fd_sc_hd__nand2_1 _06315_ (.A(\core.CPU_Dmem_value_a5[15][15] ),
    .B(net451),
    .Y(_01754_));
 sky130_fd_sc_hd__a21oi_1 _06316_ (.A1(_01753_),
    .A2(_01754_),
    .B1(net603),
    .Y(_00406_));
 sky130_fd_sc_hd__nand2_1 _06318_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net515),
    .Y(_01756_));
 sky130_fd_sc_hd__nand2_1 _06320_ (.A(\core.CPU_Dmem_value_a5[15][16] ),
    .B(net451),
    .Y(_01758_));
 sky130_fd_sc_hd__a21oi_1 _06321_ (.A1(_01756_),
    .A2(_01758_),
    .B1(net604),
    .Y(_00407_));
 sky130_fd_sc_hd__nand2_1 _06322_ (.A(net579),
    .B(net515),
    .Y(_01759_));
 sky130_fd_sc_hd__nand2_1 _06323_ (.A(\core.CPU_Dmem_value_a5[15][17] ),
    .B(net451),
    .Y(_01760_));
 sky130_fd_sc_hd__a21oi_1 _06324_ (.A1(_01759_),
    .A2(_01760_),
    .B1(net604),
    .Y(_00408_));
 sky130_fd_sc_hd__nand2_1 _06325_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net515),
    .Y(_01761_));
 sky130_fd_sc_hd__nand2_1 _06326_ (.A(\core.CPU_Dmem_value_a5[15][18] ),
    .B(net451),
    .Y(_01762_));
 sky130_fd_sc_hd__a21oi_1 _06327_ (.A1(_01761_),
    .A2(_01762_),
    .B1(net604),
    .Y(_00409_));
 sky130_fd_sc_hd__nand2_1 _06328_ (.A(net578),
    .B(net516),
    .Y(_01763_));
 sky130_fd_sc_hd__nand2_1 _06329_ (.A(\core.CPU_Dmem_value_a5[15][19] ),
    .B(_01735_),
    .Y(_01764_));
 sky130_fd_sc_hd__a21oi_1 _06330_ (.A1(_01763_),
    .A2(_01764_),
    .B1(net600),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _06331_ (.A(\core.CPU_Dmem_value_a5[15][1] ),
    .B(net451),
    .Y(_01765_));
 sky130_fd_sc_hd__nand2_1 _06332_ (.A(net577),
    .B(net515),
    .Y(_01766_));
 sky130_fd_sc_hd__nand3b_1 _06333_ (.A_N(net605),
    .B(_01765_),
    .C(_01766_),
    .Y(_00411_));
 sky130_fd_sc_hd__nand2_1 _06334_ (.A(net576),
    .B(net516),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_1 _06335_ (.A(\core.CPU_Dmem_value_a5[15][20] ),
    .B(net451),
    .Y(_01768_));
 sky130_fd_sc_hd__a21oi_1 _06336_ (.A1(_01767_),
    .A2(_01768_),
    .B1(net601),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _06337_ (.A(net575),
    .B(net516),
    .Y(_01769_));
 sky130_fd_sc_hd__nand2_1 _06338_ (.A(\core.CPU_Dmem_value_a5[15][21] ),
    .B(net451),
    .Y(_01770_));
 sky130_fd_sc_hd__a21oi_1 _06340_ (.A1(_01769_),
    .A2(_01770_),
    .B1(net601),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_1 _06341_ (.A(net574),
    .B(net516),
    .Y(_01772_));
 sky130_fd_sc_hd__nand2_1 _06342_ (.A(\core.CPU_Dmem_value_a5[15][22] ),
    .B(_01735_),
    .Y(_01773_));
 sky130_fd_sc_hd__a21oi_1 _06343_ (.A1(_01772_),
    .A2(_01773_),
    .B1(net601),
    .Y(_00414_));
 sky130_fd_sc_hd__nand2_1 _06344_ (.A(net573),
    .B(net516),
    .Y(_01774_));
 sky130_fd_sc_hd__nand2_1 _06345_ (.A(\core.CPU_Dmem_value_a5[15][23] ),
    .B(_01735_),
    .Y(_01775_));
 sky130_fd_sc_hd__a21oi_1 _06346_ (.A1(_01774_),
    .A2(_01775_),
    .B1(net601),
    .Y(_00415_));
 sky130_fd_sc_hd__nand2_1 _06347_ (.A(net572),
    .B(net516),
    .Y(_01776_));
 sky130_fd_sc_hd__nand2_1 _06348_ (.A(\core.CPU_Dmem_value_a5[15][24] ),
    .B(_01735_),
    .Y(_01777_));
 sky130_fd_sc_hd__a21oi_1 _06349_ (.A1(_01776_),
    .A2(_01777_),
    .B1(net601),
    .Y(_00416_));
 sky130_fd_sc_hd__nand2_1 _06350_ (.A(net571),
    .B(net516),
    .Y(_01778_));
 sky130_fd_sc_hd__nand2_1 _06351_ (.A(\core.CPU_Dmem_value_a5[15][25] ),
    .B(_01735_),
    .Y(_01779_));
 sky130_fd_sc_hd__a21oi_1 _06352_ (.A1(_01778_),
    .A2(_01779_),
    .B1(net601),
    .Y(_00417_));
 sky130_fd_sc_hd__nand2_1 _06354_ (.A(net570),
    .B(net515),
    .Y(_01781_));
 sky130_fd_sc_hd__nand2_1 _06356_ (.A(\core.CPU_Dmem_value_a5[15][26] ),
    .B(net451),
    .Y(_01783_));
 sky130_fd_sc_hd__a21oi_1 _06357_ (.A1(_01781_),
    .A2(_01783_),
    .B1(net603),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _06358_ (.A(net569),
    .B(net515),
    .Y(_01784_));
 sky130_fd_sc_hd__nand2_1 _06359_ (.A(\core.CPU_Dmem_value_a5[15][27] ),
    .B(net451),
    .Y(_01785_));
 sky130_fd_sc_hd__a21oi_1 _06360_ (.A1(_01784_),
    .A2(_01785_),
    .B1(net604),
    .Y(_00419_));
 sky130_fd_sc_hd__nand2_1 _06361_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net515),
    .Y(_01786_));
 sky130_fd_sc_hd__nand2_1 _06362_ (.A(\core.CPU_Dmem_value_a5[15][28] ),
    .B(net451),
    .Y(_01787_));
 sky130_fd_sc_hd__a21oi_1 _06363_ (.A1(_01786_),
    .A2(_01787_),
    .B1(net603),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _06364_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net516),
    .Y(_01788_));
 sky130_fd_sc_hd__nand2_1 _06365_ (.A(\core.CPU_Dmem_value_a5[15][29] ),
    .B(_01735_),
    .Y(_01789_));
 sky130_fd_sc_hd__a21oi_1 _06366_ (.A1(_01788_),
    .A2(_01789_),
    .B1(net599),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _06367_ (.A(\core.CPU_Dmem_value_a5[15][2] ),
    .B(net451),
    .Y(_01790_));
 sky130_fd_sc_hd__nand2_1 _06368_ (.A(net568),
    .B(net516),
    .Y(_01791_));
 sky130_fd_sc_hd__nand3b_1 _06369_ (.A_N(net605),
    .B(_01790_),
    .C(_01791_),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _06370_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net516),
    .Y(_01792_));
 sky130_fd_sc_hd__nand2_1 _06371_ (.A(\core.CPU_Dmem_value_a5[15][30] ),
    .B(_01735_),
    .Y(_01793_));
 sky130_fd_sc_hd__a21oi_1 _06372_ (.A1(_01792_),
    .A2(_01793_),
    .B1(net599),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _06373_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net516),
    .Y(_01794_));
 sky130_fd_sc_hd__nand2_1 _06374_ (.A(\core.CPU_Dmem_value_a5[15][31] ),
    .B(_01735_),
    .Y(_01795_));
 sky130_fd_sc_hd__a21oi_1 _06376_ (.A1(_01794_),
    .A2(_01795_),
    .B1(net601),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _06377_ (.A(\core.CPU_Dmem_value_a5[15][3] ),
    .B(_01735_),
    .Y(_01797_));
 sky130_fd_sc_hd__nand2_1 _06378_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net516),
    .Y(_01798_));
 sky130_fd_sc_hd__nand3b_1 _06379_ (.A_N(net599),
    .B(_01797_),
    .C(_01798_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _06380_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net515),
    .Y(_01799_));
 sky130_fd_sc_hd__nand2_1 _06381_ (.A(\core.CPU_Dmem_value_a5[15][4] ),
    .B(net451),
    .Y(_01800_));
 sky130_fd_sc_hd__a21oi_1 _06382_ (.A1(_01799_),
    .A2(_01800_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00426_));
 sky130_fd_sc_hd__nand2_1 _06383_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net515),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_1 _06384_ (.A(\core.CPU_Dmem_value_a5[15][5] ),
    .B(net451),
    .Y(_01802_));
 sky130_fd_sc_hd__a21oi_1 _06385_ (.A1(_01801_),
    .A2(_01802_),
    .B1(net605),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_1 _06386_ (.A(net567),
    .B(net516),
    .Y(_01803_));
 sky130_fd_sc_hd__nand2_1 _06387_ (.A(\core.CPU_Dmem_value_a5[15][6] ),
    .B(_01735_),
    .Y(_01804_));
 sky130_fd_sc_hd__a21oi_1 _06388_ (.A1(_01803_),
    .A2(_01804_),
    .B1(net602),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _06389_ (.A(net566),
    .B(net516),
    .Y(_01805_));
 sky130_fd_sc_hd__nand2_1 _06390_ (.A(\core.CPU_Dmem_value_a5[15][7] ),
    .B(_01735_),
    .Y(_01806_));
 sky130_fd_sc_hd__a21oi_1 _06391_ (.A1(_01805_),
    .A2(_01806_),
    .B1(net602),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _06392_ (.A(net565),
    .B(net516),
    .Y(_01807_));
 sky130_fd_sc_hd__nand2_1 _06393_ (.A(\core.CPU_Dmem_value_a5[15][8] ),
    .B(_01735_),
    .Y(_01808_));
 sky130_fd_sc_hd__a21oi_1 _06394_ (.A1(_01807_),
    .A2(_01808_),
    .B1(net601),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _06395_ (.A(net564),
    .B(net516),
    .Y(_01809_));
 sky130_fd_sc_hd__nand2_1 _06396_ (.A(\core.CPU_Dmem_value_a5[15][9] ),
    .B(net451),
    .Y(_01810_));
 sky130_fd_sc_hd__a21oi_1 _06397_ (.A1(_01809_),
    .A2(_01810_),
    .B1(net603),
    .Y(_00431_));
 sky130_fd_sc_hd__nor3_2 _06398_ (.A(\core.CPU_dmem_addr_a4[3] ),
    .B(\core.CPU_dmem_addr_a4[2] ),
    .C(_01580_),
    .Y(_01811_));
 sky130_fd_sc_hd__nand2_2 _06400_ (.A(net560),
    .B(net514),
    .Y(_01813_));
 sky130_fd_sc_hd__nand2_1 _06402_ (.A(\core.CPU_Dmem_value_a5[1][0] ),
    .B(net450),
    .Y(_01815_));
 sky130_fd_sc_hd__nor4_2 _06403_ (.A(\core.CPU_dmem_addr_a4[3] ),
    .B(\core.CPU_dmem_addr_a4[2] ),
    .C(net561),
    .D(_01580_),
    .Y(_01816_));
 sky130_fd_sc_hd__nand2_1 _06405_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net512),
    .Y(_01818_));
 sky130_fd_sc_hd__nand3b_1 _06406_ (.A_N(\core.CPU_reset_a4 ),
    .B(_01815_),
    .C(_01818_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _06407_ (.A(net584),
    .B(net511),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_1 _06408_ (.A(\core.CPU_Dmem_value_a5[1][10] ),
    .B(_01813_),
    .Y(_01820_));
 sky130_fd_sc_hd__a21oi_1 _06409_ (.A1(_01819_),
    .A2(_01820_),
    .B1(net601),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _06410_ (.A(net583),
    .B(net511),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_1 _06411_ (.A(\core.CPU_Dmem_value_a5[1][11] ),
    .B(_01813_),
    .Y(_01822_));
 sky130_fd_sc_hd__a21oi_1 _06412_ (.A1(_01821_),
    .A2(_01822_),
    .B1(net600),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _06413_ (.A(net582),
    .B(net511),
    .Y(_01823_));
 sky130_fd_sc_hd__nand2_1 _06414_ (.A(\core.CPU_Dmem_value_a5[1][12] ),
    .B(_01813_),
    .Y(_01824_));
 sky130_fd_sc_hd__a21oi_1 _06415_ (.A1(_01823_),
    .A2(_01824_),
    .B1(net602),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _06416_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net512),
    .Y(_01825_));
 sky130_fd_sc_hd__nand2_1 _06417_ (.A(\core.CPU_Dmem_value_a5[1][13] ),
    .B(net450),
    .Y(_01826_));
 sky130_fd_sc_hd__a21oi_1 _06419_ (.A1(_01825_),
    .A2(_01826_),
    .B1(net604),
    .Y(_00436_));
 sky130_fd_sc_hd__nand2_1 _06420_ (.A(net581),
    .B(net511),
    .Y(_01828_));
 sky130_fd_sc_hd__nand2_1 _06421_ (.A(\core.CPU_Dmem_value_a5[1][14] ),
    .B(net450),
    .Y(_01829_));
 sky130_fd_sc_hd__a21oi_1 _06422_ (.A1(_01828_),
    .A2(_01829_),
    .B1(net599),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _06423_ (.A(net580),
    .B(net512),
    .Y(_01830_));
 sky130_fd_sc_hd__nand2_1 _06424_ (.A(\core.CPU_Dmem_value_a5[1][15] ),
    .B(net450),
    .Y(_01831_));
 sky130_fd_sc_hd__a21oi_1 _06425_ (.A1(_01830_),
    .A2(_01831_),
    .B1(net603),
    .Y(_00438_));
 sky130_fd_sc_hd__nand2_1 _06426_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net512),
    .Y(_01832_));
 sky130_fd_sc_hd__nand2_1 _06427_ (.A(\core.CPU_Dmem_value_a5[1][16] ),
    .B(net450),
    .Y(_01833_));
 sky130_fd_sc_hd__a21oi_1 _06428_ (.A1(_01832_),
    .A2(_01833_),
    .B1(net604),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _06429_ (.A(net579),
    .B(net512),
    .Y(_01834_));
 sky130_fd_sc_hd__nand2_1 _06430_ (.A(\core.CPU_Dmem_value_a5[1][17] ),
    .B(net450),
    .Y(_01835_));
 sky130_fd_sc_hd__a21oi_1 _06431_ (.A1(_01834_),
    .A2(_01835_),
    .B1(net604),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _06432_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net512),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_1 _06433_ (.A(\core.CPU_Dmem_value_a5[1][18] ),
    .B(net450),
    .Y(_01837_));
 sky130_fd_sc_hd__a21oi_1 _06434_ (.A1(_01836_),
    .A2(_01837_),
    .B1(net604),
    .Y(_00441_));
 sky130_fd_sc_hd__nand2_1 _06436_ (.A(net578),
    .B(net511),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _06438_ (.A(\core.CPU_Dmem_value_a5[1][19] ),
    .B(net450),
    .Y(_01841_));
 sky130_fd_sc_hd__a21oi_1 _06439_ (.A1(_01839_),
    .A2(_01841_),
    .B1(net600),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_1 _06440_ (.A(net577),
    .B(net512),
    .Y(_01842_));
 sky130_fd_sc_hd__nand2_1 _06441_ (.A(\core.CPU_Dmem_value_a5[1][1] ),
    .B(net450),
    .Y(_01843_));
 sky130_fd_sc_hd__a21oi_1 _06442_ (.A1(_01842_),
    .A2(_01843_),
    .B1(net605),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_1 _06443_ (.A(net576),
    .B(net512),
    .Y(_01844_));
 sky130_fd_sc_hd__nand2_1 _06444_ (.A(\core.CPU_Dmem_value_a5[1][20] ),
    .B(net450),
    .Y(_01845_));
 sky130_fd_sc_hd__a21oi_1 _06445_ (.A1(_01844_),
    .A2(_01845_),
    .B1(net601),
    .Y(_00444_));
 sky130_fd_sc_hd__nand2_1 _06446_ (.A(net575),
    .B(net512),
    .Y(_01846_));
 sky130_fd_sc_hd__nand2_1 _06447_ (.A(\core.CPU_Dmem_value_a5[1][21] ),
    .B(net450),
    .Y(_01847_));
 sky130_fd_sc_hd__a21oi_1 _06448_ (.A1(_01846_),
    .A2(_01847_),
    .B1(net603),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2_1 _06449_ (.A(net574),
    .B(net511),
    .Y(_01848_));
 sky130_fd_sc_hd__nand2_1 _06450_ (.A(\core.CPU_Dmem_value_a5[1][22] ),
    .B(_01813_),
    .Y(_01849_));
 sky130_fd_sc_hd__a21oi_1 _06452_ (.A1(_01848_),
    .A2(_01849_),
    .B1(net601),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_1 _06453_ (.A(net573),
    .B(net511),
    .Y(_01851_));
 sky130_fd_sc_hd__nand2_1 _06454_ (.A(\core.CPU_Dmem_value_a5[1][23] ),
    .B(_01813_),
    .Y(_01852_));
 sky130_fd_sc_hd__a21oi_1 _06455_ (.A1(_01851_),
    .A2(_01852_),
    .B1(net601),
    .Y(_00447_));
 sky130_fd_sc_hd__nand2_1 _06456_ (.A(net572),
    .B(net511),
    .Y(_01853_));
 sky130_fd_sc_hd__nand2_1 _06457_ (.A(\core.CPU_Dmem_value_a5[1][24] ),
    .B(net450),
    .Y(_01854_));
 sky130_fd_sc_hd__a21oi_1 _06458_ (.A1(_01853_),
    .A2(_01854_),
    .B1(net600),
    .Y(_00448_));
 sky130_fd_sc_hd__nand2_1 _06459_ (.A(net571),
    .B(net512),
    .Y(_01855_));
 sky130_fd_sc_hd__nand2_1 _06460_ (.A(\core.CPU_Dmem_value_a5[1][25] ),
    .B(net450),
    .Y(_01856_));
 sky130_fd_sc_hd__a21oi_1 _06461_ (.A1(_01855_),
    .A2(_01856_),
    .B1(net601),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _06462_ (.A(net570),
    .B(net512),
    .Y(_01857_));
 sky130_fd_sc_hd__nand2_1 _06463_ (.A(\core.CPU_Dmem_value_a5[1][26] ),
    .B(net450),
    .Y(_01858_));
 sky130_fd_sc_hd__a21oi_1 _06464_ (.A1(_01857_),
    .A2(_01858_),
    .B1(net603),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _06465_ (.A(net569),
    .B(net512),
    .Y(_01859_));
 sky130_fd_sc_hd__nand2_1 _06466_ (.A(\core.CPU_Dmem_value_a5[1][27] ),
    .B(net450),
    .Y(_01860_));
 sky130_fd_sc_hd__a21oi_1 _06467_ (.A1(_01859_),
    .A2(_01860_),
    .B1(net604),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _06469_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net512),
    .Y(_01862_));
 sky130_fd_sc_hd__nand2_1 _06471_ (.A(\core.CPU_Dmem_value_a5[1][28] ),
    .B(net450),
    .Y(_01864_));
 sky130_fd_sc_hd__a21oi_1 _06472_ (.A1(_01862_),
    .A2(_01864_),
    .B1(net600),
    .Y(_00452_));
 sky130_fd_sc_hd__nand2_1 _06473_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net511),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _06474_ (.A(\core.CPU_Dmem_value_a5[1][29] ),
    .B(net450),
    .Y(_01866_));
 sky130_fd_sc_hd__a21oi_1 _06475_ (.A1(_01865_),
    .A2(_01866_),
    .B1(net602),
    .Y(_00453_));
 sky130_fd_sc_hd__nand2_1 _06476_ (.A(net568),
    .B(net512),
    .Y(_01867_));
 sky130_fd_sc_hd__nand2_1 _06477_ (.A(\core.CPU_Dmem_value_a5[1][2] ),
    .B(net450),
    .Y(_01868_));
 sky130_fd_sc_hd__a21oi_1 _06478_ (.A1(_01867_),
    .A2(_01868_),
    .B1(net605),
    .Y(_00454_));
 sky130_fd_sc_hd__nand2_1 _06479_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net511),
    .Y(_01869_));
 sky130_fd_sc_hd__nand2_1 _06480_ (.A(\core.CPU_Dmem_value_a5[1][30] ),
    .B(net450),
    .Y(_01870_));
 sky130_fd_sc_hd__a21oi_1 _06481_ (.A1(_01869_),
    .A2(_01870_),
    .B1(net602),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_1 _06482_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net512),
    .Y(_01871_));
 sky130_fd_sc_hd__nand2_1 _06483_ (.A(\core.CPU_Dmem_value_a5[1][31] ),
    .B(_01813_),
    .Y(_01872_));
 sky130_fd_sc_hd__a21oi_1 _06485_ (.A1(_01871_),
    .A2(_01872_),
    .B1(net601),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _06486_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net511),
    .Y(_01874_));
 sky130_fd_sc_hd__nand2_1 _06487_ (.A(\core.CPU_Dmem_value_a5[1][3] ),
    .B(net450),
    .Y(_01875_));
 sky130_fd_sc_hd__a21oi_1 _06488_ (.A1(_01874_),
    .A2(_01875_),
    .B1(net599),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_1 _06489_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net512),
    .Y(_01876_));
 sky130_fd_sc_hd__nand2_1 _06490_ (.A(\core.CPU_Dmem_value_a5[1][4] ),
    .B(net450),
    .Y(_01877_));
 sky130_fd_sc_hd__a21oi_1 _06491_ (.A1(_01876_),
    .A2(_01877_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _06492_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net512),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _06493_ (.A(\core.CPU_Dmem_value_a5[1][5] ),
    .B(net450),
    .Y(_01879_));
 sky130_fd_sc_hd__a21oi_1 _06494_ (.A1(_01878_),
    .A2(_01879_),
    .B1(net605),
    .Y(_00459_));
 sky130_fd_sc_hd__nand2_1 _06495_ (.A(net567),
    .B(net511),
    .Y(_01880_));
 sky130_fd_sc_hd__nand2_1 _06496_ (.A(\core.CPU_Dmem_value_a5[1][6] ),
    .B(net450),
    .Y(_01881_));
 sky130_fd_sc_hd__a21oi_1 _06497_ (.A1(_01880_),
    .A2(_01881_),
    .B1(net599),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2_1 _06498_ (.A(net566),
    .B(net511),
    .Y(_01882_));
 sky130_fd_sc_hd__nand2_1 _06499_ (.A(\core.CPU_Dmem_value_a5[1][7] ),
    .B(net450),
    .Y(_01883_));
 sky130_fd_sc_hd__a21oi_1 _06500_ (.A1(_01882_),
    .A2(_01883_),
    .B1(net599),
    .Y(_00461_));
 sky130_fd_sc_hd__nand2_1 _06501_ (.A(net565),
    .B(net512),
    .Y(_01884_));
 sky130_fd_sc_hd__nand2_1 _06502_ (.A(\core.CPU_Dmem_value_a5[1][8] ),
    .B(_01813_),
    .Y(_01885_));
 sky130_fd_sc_hd__a21oi_1 _06503_ (.A1(_01884_),
    .A2(_01885_),
    .B1(net601),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _06504_ (.A(net564),
    .B(net512),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_1 _06505_ (.A(\core.CPU_Dmem_value_a5[1][9] ),
    .B(net450),
    .Y(_01887_));
 sky130_fd_sc_hd__a21oi_1 _06506_ (.A1(_01886_),
    .A2(_01887_),
    .B1(net605),
    .Y(_00463_));
 sky130_fd_sc_hd__nor4_2 _06507_ (.A(\core.CPU_dmem_addr_a4[3] ),
    .B(\core.CPU_dmem_addr_a4[2] ),
    .C(net561),
    .D(_01344_),
    .Y(_01888_));
 sky130_fd_sc_hd__nand2_1 _06509_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net509),
    .Y(_01890_));
 sky130_fd_sc_hd__nor3_2 _06510_ (.A(\core.CPU_dmem_addr_a4[3] ),
    .B(\core.CPU_dmem_addr_a4[2] ),
    .C(_01344_),
    .Y(_01891_));
 sky130_fd_sc_hd__nand2_2 _06512_ (.A(net560),
    .B(net508),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2_1 _06514_ (.A(\core.CPU_Dmem_value_a5[2][0] ),
    .B(net449),
    .Y(_01895_));
 sky130_fd_sc_hd__a21oi_1 _06515_ (.A1(_01890_),
    .A2(_01895_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00464_));
 sky130_fd_sc_hd__nand2_1 _06516_ (.A(net584),
    .B(net510),
    .Y(_01896_));
 sky130_fd_sc_hd__nand2_1 _06517_ (.A(\core.CPU_Dmem_value_a5[2][10] ),
    .B(net449),
    .Y(_01897_));
 sky130_fd_sc_hd__a21oi_1 _06518_ (.A1(_01896_),
    .A2(_01897_),
    .B1(net601),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _06519_ (.A(net583),
    .B(net510),
    .Y(_01898_));
 sky130_fd_sc_hd__nand2_1 _06520_ (.A(\core.CPU_Dmem_value_a5[2][11] ),
    .B(net449),
    .Y(_01899_));
 sky130_fd_sc_hd__a21oi_1 _06522_ (.A1(_01898_),
    .A2(_01899_),
    .B1(net600),
    .Y(_00466_));
 sky130_fd_sc_hd__nand2_1 _06523_ (.A(net582),
    .B(net510),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2_1 _06524_ (.A(\core.CPU_Dmem_value_a5[2][12] ),
    .B(net449),
    .Y(_01902_));
 sky130_fd_sc_hd__a21oi_1 _06525_ (.A1(_01901_),
    .A2(_01902_),
    .B1(net602),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _06526_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net509),
    .Y(_01903_));
 sky130_fd_sc_hd__nand2_1 _06527_ (.A(\core.CPU_Dmem_value_a5[2][13] ),
    .B(net449),
    .Y(_01904_));
 sky130_fd_sc_hd__a21oi_1 _06528_ (.A1(_01903_),
    .A2(_01904_),
    .B1(net604),
    .Y(_00468_));
 sky130_fd_sc_hd__nand2_1 _06529_ (.A(net581),
    .B(net510),
    .Y(_01905_));
 sky130_fd_sc_hd__nand2_1 _06530_ (.A(\core.CPU_Dmem_value_a5[2][14] ),
    .B(_01893_),
    .Y(_01906_));
 sky130_fd_sc_hd__a21oi_1 _06531_ (.A1(_01905_),
    .A2(_01906_),
    .B1(net599),
    .Y(_00469_));
 sky130_fd_sc_hd__nand2_1 _06532_ (.A(net580),
    .B(net510),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _06533_ (.A(\core.CPU_Dmem_value_a5[2][15] ),
    .B(net449),
    .Y(_01908_));
 sky130_fd_sc_hd__a21oi_1 _06534_ (.A1(_01907_),
    .A2(_01908_),
    .B1(net601),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _06535_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net509),
    .Y(_01909_));
 sky130_fd_sc_hd__nand2_1 _06536_ (.A(\core.CPU_Dmem_value_a5[2][16] ),
    .B(net449),
    .Y(_01910_));
 sky130_fd_sc_hd__a21oi_1 _06537_ (.A1(_01909_),
    .A2(_01910_),
    .B1(net604),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _06538_ (.A(net579),
    .B(net509),
    .Y(_01911_));
 sky130_fd_sc_hd__nand2_1 _06539_ (.A(\core.CPU_Dmem_value_a5[2][17] ),
    .B(net449),
    .Y(_01912_));
 sky130_fd_sc_hd__a21oi_1 _06540_ (.A1(_01911_),
    .A2(_01912_),
    .B1(net604),
    .Y(_00472_));
 sky130_fd_sc_hd__nand2_1 _06542_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net509),
    .Y(_01914_));
 sky130_fd_sc_hd__nand2_1 _06544_ (.A(\core.CPU_Dmem_value_a5[2][18] ),
    .B(net449),
    .Y(_01916_));
 sky130_fd_sc_hd__a21oi_1 _06545_ (.A1(_01914_),
    .A2(_01916_),
    .B1(net604),
    .Y(_00473_));
 sky130_fd_sc_hd__nand2_1 _06546_ (.A(net578),
    .B(net510),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_1 _06547_ (.A(\core.CPU_Dmem_value_a5[2][19] ),
    .B(_01893_),
    .Y(_01918_));
 sky130_fd_sc_hd__a21oi_1 _06548_ (.A1(_01917_),
    .A2(_01918_),
    .B1(net600),
    .Y(_00474_));
 sky130_fd_sc_hd__nand2_1 _06549_ (.A(\core.CPU_Dmem_value_a5[2][1] ),
    .B(net449),
    .Y(_01919_));
 sky130_fd_sc_hd__nand2_1 _06550_ (.A(net577),
    .B(net510),
    .Y(_01920_));
 sky130_fd_sc_hd__nand3b_1 _06551_ (.A_N(net605),
    .B(_01919_),
    .C(_01920_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_1 _06552_ (.A(net576),
    .B(net510),
    .Y(_01921_));
 sky130_fd_sc_hd__nand2_1 _06553_ (.A(\core.CPU_Dmem_value_a5[2][20] ),
    .B(net449),
    .Y(_01922_));
 sky130_fd_sc_hd__a21oi_1 _06554_ (.A1(_01921_),
    .A2(_01922_),
    .B1(net601),
    .Y(_00476_));
 sky130_fd_sc_hd__nand2_1 _06555_ (.A(net575),
    .B(net510),
    .Y(_01923_));
 sky130_fd_sc_hd__nand2_1 _06556_ (.A(\core.CPU_Dmem_value_a5[2][21] ),
    .B(net449),
    .Y(_01924_));
 sky130_fd_sc_hd__a21oi_1 _06558_ (.A1(_01923_),
    .A2(_01924_),
    .B1(net603),
    .Y(_00477_));
 sky130_fd_sc_hd__nand2_1 _06559_ (.A(net574),
    .B(net510),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_1 _06560_ (.A(\core.CPU_Dmem_value_a5[2][22] ),
    .B(net449),
    .Y(_01927_));
 sky130_fd_sc_hd__a21oi_1 _06561_ (.A1(_01926_),
    .A2(_01927_),
    .B1(net601),
    .Y(_00478_));
 sky130_fd_sc_hd__nand2_1 _06562_ (.A(net573),
    .B(net510),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _06563_ (.A(\core.CPU_Dmem_value_a5[2][23] ),
    .B(net449),
    .Y(_01929_));
 sky130_fd_sc_hd__a21oi_1 _06564_ (.A1(_01928_),
    .A2(_01929_),
    .B1(net601),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _06565_ (.A(net572),
    .B(net510),
    .Y(_01930_));
 sky130_fd_sc_hd__nand2_1 _06566_ (.A(\core.CPU_Dmem_value_a5[2][24] ),
    .B(net449),
    .Y(_01931_));
 sky130_fd_sc_hd__a21oi_1 _06567_ (.A1(_01930_),
    .A2(_01931_),
    .B1(net601),
    .Y(_00480_));
 sky130_fd_sc_hd__nand2_1 _06568_ (.A(net571),
    .B(net510),
    .Y(_01932_));
 sky130_fd_sc_hd__nand2_1 _06569_ (.A(\core.CPU_Dmem_value_a5[2][25] ),
    .B(_01893_),
    .Y(_01933_));
 sky130_fd_sc_hd__a21oi_1 _06570_ (.A1(_01932_),
    .A2(_01933_),
    .B1(net601),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _06571_ (.A(net570),
    .B(net510),
    .Y(_01934_));
 sky130_fd_sc_hd__nand2_1 _06572_ (.A(\core.CPU_Dmem_value_a5[2][26] ),
    .B(net449),
    .Y(_01935_));
 sky130_fd_sc_hd__a21oi_1 _06573_ (.A1(_01934_),
    .A2(_01935_),
    .B1(net603),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _06574_ (.A(net569),
    .B(net509),
    .Y(_01936_));
 sky130_fd_sc_hd__nand2_1 _06575_ (.A(\core.CPU_Dmem_value_a5[2][27] ),
    .B(net449),
    .Y(_01937_));
 sky130_fd_sc_hd__a21oi_1 _06576_ (.A1(_01936_),
    .A2(_01937_),
    .B1(net604),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _06578_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net510),
    .Y(_01939_));
 sky130_fd_sc_hd__nand2_1 _06580_ (.A(\core.CPU_Dmem_value_a5[2][28] ),
    .B(net449),
    .Y(_01941_));
 sky130_fd_sc_hd__a21oi_1 _06581_ (.A1(_01939_),
    .A2(_01941_),
    .B1(net603),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _06582_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net510),
    .Y(_01942_));
 sky130_fd_sc_hd__nand2_1 _06583_ (.A(\core.CPU_Dmem_value_a5[2][29] ),
    .B(_01893_),
    .Y(_01943_));
 sky130_fd_sc_hd__a21oi_1 _06584_ (.A1(_01942_),
    .A2(_01943_),
    .B1(net599),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_1 _06585_ (.A(net568),
    .B(net510),
    .Y(_01944_));
 sky130_fd_sc_hd__nand2_1 _06586_ (.A(\core.CPU_Dmem_value_a5[2][2] ),
    .B(net449),
    .Y(_01945_));
 sky130_fd_sc_hd__a21oi_1 _06587_ (.A1(_01944_),
    .A2(_01945_),
    .B1(net605),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _06588_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net510),
    .Y(_01946_));
 sky130_fd_sc_hd__nand2_1 _06589_ (.A(\core.CPU_Dmem_value_a5[2][30] ),
    .B(_01893_),
    .Y(_01947_));
 sky130_fd_sc_hd__a21oi_1 _06591_ (.A1(_01946_),
    .A2(_01947_),
    .B1(net602),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _06592_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net510),
    .Y(_01949_));
 sky130_fd_sc_hd__nand2_1 _06593_ (.A(\core.CPU_Dmem_value_a5[2][31] ),
    .B(net449),
    .Y(_01950_));
 sky130_fd_sc_hd__a21oi_1 _06594_ (.A1(_01949_),
    .A2(_01950_),
    .B1(net601),
    .Y(_00488_));
 sky130_fd_sc_hd__nand2_1 _06595_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net509),
    .Y(_01951_));
 sky130_fd_sc_hd__nand2_1 _06596_ (.A(\core.CPU_Dmem_value_a5[2][3] ),
    .B(net449),
    .Y(_01952_));
 sky130_fd_sc_hd__a21oi_1 _06597_ (.A1(_01951_),
    .A2(_01952_),
    .B1(net599),
    .Y(_00489_));
 sky130_fd_sc_hd__nand2_1 _06598_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net509),
    .Y(_01953_));
 sky130_fd_sc_hd__nand2_1 _06599_ (.A(\core.CPU_Dmem_value_a5[2][4] ),
    .B(net449),
    .Y(_01954_));
 sky130_fd_sc_hd__a21oi_1 _06600_ (.A1(_01953_),
    .A2(_01954_),
    .B1(net599),
    .Y(_00490_));
 sky130_fd_sc_hd__nand2_1 _06601_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net509),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _06602_ (.A(\core.CPU_Dmem_value_a5[2][5] ),
    .B(net449),
    .Y(_01956_));
 sky130_fd_sc_hd__a21oi_1 _06603_ (.A1(_01955_),
    .A2(_01956_),
    .B1(net604),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_1 _06604_ (.A(net567),
    .B(net510),
    .Y(_01957_));
 sky130_fd_sc_hd__nand2_1 _06605_ (.A(\core.CPU_Dmem_value_a5[2][6] ),
    .B(net449),
    .Y(_01958_));
 sky130_fd_sc_hd__a21oi_1 _06606_ (.A1(_01957_),
    .A2(_01958_),
    .B1(net599),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _06607_ (.A(net566),
    .B(net510),
    .Y(_01959_));
 sky130_fd_sc_hd__nand2_1 _06608_ (.A(\core.CPU_Dmem_value_a5[2][7] ),
    .B(net449),
    .Y(_01960_));
 sky130_fd_sc_hd__a21oi_1 _06609_ (.A1(_01959_),
    .A2(_01960_),
    .B1(net602),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _06610_ (.A(net565),
    .B(net510),
    .Y(_01961_));
 sky130_fd_sc_hd__nand2_1 _06611_ (.A(\core.CPU_Dmem_value_a5[2][8] ),
    .B(net449),
    .Y(_01962_));
 sky130_fd_sc_hd__a21oi_1 _06612_ (.A1(_01961_),
    .A2(_01962_),
    .B1(net601),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _06613_ (.A(net564),
    .B(net510),
    .Y(_01963_));
 sky130_fd_sc_hd__nand2_1 _06614_ (.A(\core.CPU_Dmem_value_a5[2][9] ),
    .B(net449),
    .Y(_01964_));
 sky130_fd_sc_hd__a21oi_1 _06615_ (.A1(_01963_),
    .A2(_01964_),
    .B1(net605),
    .Y(_00495_));
 sky130_fd_sc_hd__nor3_2 _06616_ (.A(\core.CPU_dmem_addr_a4[3] ),
    .B(\core.CPU_dmem_addr_a4[2] ),
    .C(_01425_),
    .Y(_01965_));
 sky130_fd_sc_hd__nand2_2 _06618_ (.A(net560),
    .B(net505),
    .Y(_01967_));
 sky130_fd_sc_hd__nand2_1 _06620_ (.A(\core.CPU_Dmem_value_a5[3][0] ),
    .B(net448),
    .Y(_01969_));
 sky130_fd_sc_hd__nor4_2 _06621_ (.A(\core.CPU_dmem_addr_a4[3] ),
    .B(\core.CPU_dmem_addr_a4[2] ),
    .C(net561),
    .D(_01425_),
    .Y(_01970_));
 sky130_fd_sc_hd__nand2_1 _06623_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net504),
    .Y(_01972_));
 sky130_fd_sc_hd__nand3b_1 _06624_ (.A_N(\core.CPU_reset_a4 ),
    .B(_01969_),
    .C(_01972_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _06625_ (.A(net584),
    .B(net503),
    .Y(_01973_));
 sky130_fd_sc_hd__nand2_1 _06626_ (.A(\core.CPU_Dmem_value_a5[3][10] ),
    .B(net448),
    .Y(_01974_));
 sky130_fd_sc_hd__a21oi_1 _06627_ (.A1(_01973_),
    .A2(_01974_),
    .B1(net601),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _06628_ (.A(net583),
    .B(net503),
    .Y(_01975_));
 sky130_fd_sc_hd__nand2_1 _06629_ (.A(\core.CPU_Dmem_value_a5[3][11] ),
    .B(net448),
    .Y(_01976_));
 sky130_fd_sc_hd__a21oi_1 _06631_ (.A1(_01975_),
    .A2(_01976_),
    .B1(net600),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _06632_ (.A(net582),
    .B(net503),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _06633_ (.A(\core.CPU_Dmem_value_a5[3][12] ),
    .B(net448),
    .Y(_01979_));
 sky130_fd_sc_hd__a21oi_1 _06634_ (.A1(_01978_),
    .A2(_01979_),
    .B1(net602),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _06635_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net504),
    .Y(_01980_));
 sky130_fd_sc_hd__nand2_1 _06636_ (.A(\core.CPU_Dmem_value_a5[3][13] ),
    .B(net448),
    .Y(_01981_));
 sky130_fd_sc_hd__a21oi_1 _06637_ (.A1(_01980_),
    .A2(_01981_),
    .B1(net605),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_1 _06638_ (.A(net581),
    .B(net503),
    .Y(_01982_));
 sky130_fd_sc_hd__nand2_1 _06639_ (.A(\core.CPU_Dmem_value_a5[3][14] ),
    .B(_01967_),
    .Y(_01983_));
 sky130_fd_sc_hd__a21oi_1 _06640_ (.A1(_01982_),
    .A2(_01983_),
    .B1(net602),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _06641_ (.A(net580),
    .B(net504),
    .Y(_01984_));
 sky130_fd_sc_hd__nand2_1 _06642_ (.A(\core.CPU_Dmem_value_a5[3][15] ),
    .B(net448),
    .Y(_01985_));
 sky130_fd_sc_hd__a21oi_1 _06643_ (.A1(_01984_),
    .A2(_01985_),
    .B1(net603),
    .Y(_00502_));
 sky130_fd_sc_hd__nand2_1 _06644_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net504),
    .Y(_01986_));
 sky130_fd_sc_hd__nand2_1 _06645_ (.A(\core.CPU_Dmem_value_a5[3][16] ),
    .B(net448),
    .Y(_01987_));
 sky130_fd_sc_hd__a21oi_1 _06646_ (.A1(_01986_),
    .A2(_01987_),
    .B1(net604),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _06647_ (.A(net579),
    .B(net504),
    .Y(_01988_));
 sky130_fd_sc_hd__nand2_1 _06648_ (.A(\core.CPU_Dmem_value_a5[3][17] ),
    .B(net448),
    .Y(_01989_));
 sky130_fd_sc_hd__a21oi_1 _06649_ (.A1(_01988_),
    .A2(_01989_),
    .B1(net604),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _06651_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net504),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_1 _06653_ (.A(\core.CPU_Dmem_value_a5[3][18] ),
    .B(net448),
    .Y(_01993_));
 sky130_fd_sc_hd__a21oi_1 _06654_ (.A1(_01991_),
    .A2(_01993_),
    .B1(net604),
    .Y(_00505_));
 sky130_fd_sc_hd__nand2_1 _06655_ (.A(net578),
    .B(net503),
    .Y(_01994_));
 sky130_fd_sc_hd__nand2_1 _06656_ (.A(\core.CPU_Dmem_value_a5[3][19] ),
    .B(_01967_),
    .Y(_01995_));
 sky130_fd_sc_hd__a21oi_1 _06657_ (.A1(_01994_),
    .A2(_01995_),
    .B1(net600),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _06659_ (.A(\core.CPU_Dmem_value_a5[3][1] ),
    .B(net448),
    .Y(_01997_));
 sky130_fd_sc_hd__nand2_1 _06660_ (.A(net577),
    .B(net504),
    .Y(_01998_));
 sky130_fd_sc_hd__nand3b_1 _06661_ (.A_N(net605),
    .B(_01997_),
    .C(_01998_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _06662_ (.A(net576),
    .B(net503),
    .Y(_01999_));
 sky130_fd_sc_hd__nand2_1 _06663_ (.A(\core.CPU_Dmem_value_a5[3][20] ),
    .B(net448),
    .Y(_02000_));
 sky130_fd_sc_hd__a21oi_1 _06664_ (.A1(_01999_),
    .A2(_02000_),
    .B1(net601),
    .Y(_00508_));
 sky130_fd_sc_hd__nand2_1 _06665_ (.A(net575),
    .B(net504),
    .Y(_02001_));
 sky130_fd_sc_hd__nand2_1 _06666_ (.A(\core.CPU_Dmem_value_a5[3][21] ),
    .B(net448),
    .Y(_02002_));
 sky130_fd_sc_hd__a21oi_1 _06669_ (.A1(_02001_),
    .A2(_02002_),
    .B1(net605),
    .Y(_00509_));
 sky130_fd_sc_hd__nand2_1 _06670_ (.A(net574),
    .B(net503),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _06671_ (.A(\core.CPU_Dmem_value_a5[3][22] ),
    .B(net448),
    .Y(_02006_));
 sky130_fd_sc_hd__a21oi_1 _06672_ (.A1(_02005_),
    .A2(_02006_),
    .B1(net601),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _06673_ (.A(net573),
    .B(net503),
    .Y(_02007_));
 sky130_fd_sc_hd__nand2_1 _06674_ (.A(\core.CPU_Dmem_value_a5[3][23] ),
    .B(net448),
    .Y(_02008_));
 sky130_fd_sc_hd__a21oi_1 _06675_ (.A1(_02007_),
    .A2(_02008_),
    .B1(net601),
    .Y(_00511_));
 sky130_fd_sc_hd__nand2_1 _06676_ (.A(net572),
    .B(net503),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_1 _06677_ (.A(\core.CPU_Dmem_value_a5[3][24] ),
    .B(net448),
    .Y(_02010_));
 sky130_fd_sc_hd__a21oi_1 _06678_ (.A1(_02009_),
    .A2(_02010_),
    .B1(net601),
    .Y(_00512_));
 sky130_fd_sc_hd__nand2_1 _06679_ (.A(net571),
    .B(net503),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2_1 _06680_ (.A(\core.CPU_Dmem_value_a5[3][25] ),
    .B(_01967_),
    .Y(_02012_));
 sky130_fd_sc_hd__a21oi_1 _06681_ (.A1(_02011_),
    .A2(_02012_),
    .B1(net601),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _06682_ (.A(net570),
    .B(net504),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_1 _06683_ (.A(\core.CPU_Dmem_value_a5[3][26] ),
    .B(net448),
    .Y(_02014_));
 sky130_fd_sc_hd__a21oi_1 _06684_ (.A1(_02013_),
    .A2(_02014_),
    .B1(net603),
    .Y(_00514_));
 sky130_fd_sc_hd__nand2_1 _06685_ (.A(net569),
    .B(net504),
    .Y(_02015_));
 sky130_fd_sc_hd__nand2_1 _06686_ (.A(\core.CPU_Dmem_value_a5[3][27] ),
    .B(net448),
    .Y(_02016_));
 sky130_fd_sc_hd__a21oi_1 _06687_ (.A1(_02015_),
    .A2(_02016_),
    .B1(net604),
    .Y(_00515_));
 sky130_fd_sc_hd__nand2_1 _06689_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net504),
    .Y(_02018_));
 sky130_fd_sc_hd__nand2_1 _06691_ (.A(\core.CPU_Dmem_value_a5[3][28] ),
    .B(net448),
    .Y(_02020_));
 sky130_fd_sc_hd__a21oi_1 _06692_ (.A1(_02018_),
    .A2(_02020_),
    .B1(net603),
    .Y(_00516_));
 sky130_fd_sc_hd__nand2_1 _06693_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net503),
    .Y(_02021_));
 sky130_fd_sc_hd__nand2_1 _06694_ (.A(\core.CPU_Dmem_value_a5[3][29] ),
    .B(_01967_),
    .Y(_02022_));
 sky130_fd_sc_hd__a21oi_1 _06695_ (.A1(_02021_),
    .A2(_02022_),
    .B1(net602),
    .Y(_00517_));
 sky130_fd_sc_hd__nand2_1 _06696_ (.A(net568),
    .B(net504),
    .Y(_02023_));
 sky130_fd_sc_hd__nand2_1 _06697_ (.A(\core.CPU_Dmem_value_a5[3][2] ),
    .B(net448),
    .Y(_02024_));
 sky130_fd_sc_hd__a21oi_1 _06698_ (.A1(_02023_),
    .A2(_02024_),
    .B1(net605),
    .Y(_00518_));
 sky130_fd_sc_hd__nand2_1 _06699_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net503),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_1 _06700_ (.A(\core.CPU_Dmem_value_a5[3][30] ),
    .B(_01967_),
    .Y(_02026_));
 sky130_fd_sc_hd__a21oi_1 _06702_ (.A1(_02025_),
    .A2(_02026_),
    .B1(net602),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _06703_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net504),
    .Y(_02028_));
 sky130_fd_sc_hd__nand2_1 _06704_ (.A(\core.CPU_Dmem_value_a5[3][31] ),
    .B(net448),
    .Y(_02029_));
 sky130_fd_sc_hd__a21oi_1 _06705_ (.A1(_02028_),
    .A2(_02029_),
    .B1(net601),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2_1 _06706_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(_01970_),
    .Y(_02030_));
 sky130_fd_sc_hd__nand2_1 _06707_ (.A(\core.CPU_Dmem_value_a5[3][3] ),
    .B(_01967_),
    .Y(_02031_));
 sky130_fd_sc_hd__a21oi_1 _06708_ (.A1(_02030_),
    .A2(_02031_),
    .B1(net599),
    .Y(_00521_));
 sky130_fd_sc_hd__nand2_1 _06709_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(_01970_),
    .Y(_02032_));
 sky130_fd_sc_hd__nand2_1 _06710_ (.A(\core.CPU_Dmem_value_a5[3][4] ),
    .B(_01967_),
    .Y(_02033_));
 sky130_fd_sc_hd__a21oi_1 _06711_ (.A1(_02032_),
    .A2(_02033_),
    .B1(net599),
    .Y(_00522_));
 sky130_fd_sc_hd__nand2_1 _06712_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net504),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _06713_ (.A(\core.CPU_Dmem_value_a5[3][5] ),
    .B(net448),
    .Y(_02035_));
 sky130_fd_sc_hd__a21oi_1 _06714_ (.A1(_02034_),
    .A2(_02035_),
    .B1(net605),
    .Y(_00523_));
 sky130_fd_sc_hd__nand2_1 _06715_ (.A(net567),
    .B(net503),
    .Y(_02036_));
 sky130_fd_sc_hd__nand2_1 _06716_ (.A(\core.CPU_Dmem_value_a5[3][6] ),
    .B(_01967_),
    .Y(_02037_));
 sky130_fd_sc_hd__a21oi_1 _06717_ (.A1(_02036_),
    .A2(_02037_),
    .B1(net599),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_1 _06718_ (.A(net566),
    .B(net503),
    .Y(_02038_));
 sky130_fd_sc_hd__nand2_1 _06719_ (.A(\core.CPU_Dmem_value_a5[3][7] ),
    .B(_01967_),
    .Y(_02039_));
 sky130_fd_sc_hd__a21oi_1 _06720_ (.A1(_02038_),
    .A2(_02039_),
    .B1(net599),
    .Y(_00525_));
 sky130_fd_sc_hd__nand2_1 _06721_ (.A(net565),
    .B(net503),
    .Y(_02040_));
 sky130_fd_sc_hd__nand2_1 _06722_ (.A(\core.CPU_Dmem_value_a5[3][8] ),
    .B(net448),
    .Y(_02041_));
 sky130_fd_sc_hd__a21oi_1 _06723_ (.A1(_02040_),
    .A2(_02041_),
    .B1(net601),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_1 _06724_ (.A(net564),
    .B(net504),
    .Y(_02042_));
 sky130_fd_sc_hd__nand2_1 _06725_ (.A(\core.CPU_Dmem_value_a5[3][9] ),
    .B(net448),
    .Y(_02043_));
 sky130_fd_sc_hd__a21oi_1 _06726_ (.A1(_02042_),
    .A2(_02043_),
    .B1(net603),
    .Y(_00527_));
 sky130_fd_sc_hd__nand2b_1 _06727_ (.A_N(\core.CPU_dmem_addr_a4[3] ),
    .B(\core.CPU_dmem_addr_a4[2] ),
    .Y(_02044_));
 sky130_fd_sc_hd__nor4_2 _06729_ (.A(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .C(net561),
    .D(_02044_),
    .Y(_02046_));
 sky130_fd_sc_hd__nand2_1 _06731_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net501),
    .Y(_02048_));
 sky130_fd_sc_hd__nor3_2 _06732_ (.A(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .C(_02044_),
    .Y(_02049_));
 sky130_fd_sc_hd__nand2_2 _06733_ (.A(net560),
    .B(net499),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_1 _06735_ (.A(\core.CPU_Dmem_value_a5[4][0] ),
    .B(_02050_),
    .Y(_02052_));
 sky130_fd_sc_hd__a21oi_1 _06736_ (.A1(_02048_),
    .A2(_02052_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00528_));
 sky130_fd_sc_hd__nand2_1 _06737_ (.A(net584),
    .B(net502),
    .Y(_02053_));
 sky130_fd_sc_hd__nand2_1 _06738_ (.A(\core.CPU_Dmem_value_a5[4][10] ),
    .B(net447),
    .Y(_02054_));
 sky130_fd_sc_hd__a21oi_1 _06740_ (.A1(_02053_),
    .A2(_02054_),
    .B1(net601),
    .Y(_00529_));
 sky130_fd_sc_hd__nand2_1 _06741_ (.A(net583),
    .B(net502),
    .Y(_02056_));
 sky130_fd_sc_hd__nand2_1 _06742_ (.A(\core.CPU_Dmem_value_a5[4][11] ),
    .B(net447),
    .Y(_02057_));
 sky130_fd_sc_hd__a21oi_1 _06743_ (.A1(_02056_),
    .A2(_02057_),
    .B1(net600),
    .Y(_00530_));
 sky130_fd_sc_hd__nand2_1 _06744_ (.A(net582),
    .B(net502),
    .Y(_02058_));
 sky130_fd_sc_hd__nand2_1 _06745_ (.A(\core.CPU_Dmem_value_a5[4][12] ),
    .B(net447),
    .Y(_02059_));
 sky130_fd_sc_hd__a21oi_1 _06746_ (.A1(_02058_),
    .A2(_02059_),
    .B1(net602),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _06747_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net501),
    .Y(_02060_));
 sky130_fd_sc_hd__nand2_1 _06748_ (.A(\core.CPU_Dmem_value_a5[4][13] ),
    .B(net447),
    .Y(_02061_));
 sky130_fd_sc_hd__a21oi_1 _06749_ (.A1(_02060_),
    .A2(_02061_),
    .B1(net604),
    .Y(_00532_));
 sky130_fd_sc_hd__nand2_1 _06750_ (.A(net581),
    .B(net502),
    .Y(_02062_));
 sky130_fd_sc_hd__nand2_1 _06751_ (.A(\core.CPU_Dmem_value_a5[4][14] ),
    .B(_02050_),
    .Y(_02063_));
 sky130_fd_sc_hd__a21oi_1 _06752_ (.A1(_02062_),
    .A2(_02063_),
    .B1(net599),
    .Y(_00533_));
 sky130_fd_sc_hd__nand2_1 _06753_ (.A(net580),
    .B(net501),
    .Y(_02064_));
 sky130_fd_sc_hd__nand2_1 _06754_ (.A(\core.CPU_Dmem_value_a5[4][15] ),
    .B(net447),
    .Y(_02065_));
 sky130_fd_sc_hd__a21oi_1 _06755_ (.A1(_02064_),
    .A2(_02065_),
    .B1(net603),
    .Y(_00534_));
 sky130_fd_sc_hd__nand2_1 _06756_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net501),
    .Y(_02066_));
 sky130_fd_sc_hd__nand2_1 _06757_ (.A(\core.CPU_Dmem_value_a5[4][16] ),
    .B(_02050_),
    .Y(_02067_));
 sky130_fd_sc_hd__a21oi_1 _06758_ (.A1(_02066_),
    .A2(_02067_),
    .B1(net605),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _06759_ (.A(net579),
    .B(net501),
    .Y(_02068_));
 sky130_fd_sc_hd__nand2_1 _06760_ (.A(\core.CPU_Dmem_value_a5[4][17] ),
    .B(_02050_),
    .Y(_02069_));
 sky130_fd_sc_hd__a21oi_1 _06761_ (.A1(_02068_),
    .A2(_02069_),
    .B1(net604),
    .Y(_00536_));
 sky130_fd_sc_hd__nand2_1 _06763_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net501),
    .Y(_02071_));
 sky130_fd_sc_hd__nand2_1 _06765_ (.A(\core.CPU_Dmem_value_a5[4][18] ),
    .B(_02050_),
    .Y(_02073_));
 sky130_fd_sc_hd__a21oi_1 _06766_ (.A1(_02071_),
    .A2(_02073_),
    .B1(net604),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_1 _06767_ (.A(net578),
    .B(net502),
    .Y(_02074_));
 sky130_fd_sc_hd__nand2_1 _06768_ (.A(\core.CPU_Dmem_value_a5[4][19] ),
    .B(_02050_),
    .Y(_02075_));
 sky130_fd_sc_hd__a21oi_1 _06769_ (.A1(_02074_),
    .A2(_02075_),
    .B1(net600),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _06770_ (.A(net577),
    .B(net501),
    .Y(_02076_));
 sky130_fd_sc_hd__nand2_1 _06771_ (.A(\core.CPU_Dmem_value_a5[4][1] ),
    .B(net447),
    .Y(_02077_));
 sky130_fd_sc_hd__a21oi_1 _06773_ (.A1(_02076_),
    .A2(_02077_),
    .B1(net605),
    .Y(_00539_));
 sky130_fd_sc_hd__nand2_1 _06774_ (.A(net576),
    .B(net502),
    .Y(_02079_));
 sky130_fd_sc_hd__nand2_1 _06775_ (.A(\core.CPU_Dmem_value_a5[4][20] ),
    .B(net447),
    .Y(_02080_));
 sky130_fd_sc_hd__a21oi_1 _06776_ (.A1(_02079_),
    .A2(_02080_),
    .B1(net601),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_1 _06777_ (.A(net575),
    .B(net501),
    .Y(_02081_));
 sky130_fd_sc_hd__nand2_1 _06778_ (.A(\core.CPU_Dmem_value_a5[4][21] ),
    .B(net447),
    .Y(_02082_));
 sky130_fd_sc_hd__a21oi_1 _06779_ (.A1(_02081_),
    .A2(_02082_),
    .B1(net601),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_1 _06780_ (.A(net574),
    .B(net502),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _06781_ (.A(\core.CPU_Dmem_value_a5[4][22] ),
    .B(net447),
    .Y(_02084_));
 sky130_fd_sc_hd__a21oi_1 _06782_ (.A1(_02083_),
    .A2(_02084_),
    .B1(net601),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_1 _06783_ (.A(net573),
    .B(net502),
    .Y(_02085_));
 sky130_fd_sc_hd__nand2_1 _06784_ (.A(\core.CPU_Dmem_value_a5[4][23] ),
    .B(net447),
    .Y(_02086_));
 sky130_fd_sc_hd__a21oi_1 _06785_ (.A1(_02085_),
    .A2(_02086_),
    .B1(net601),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2_1 _06786_ (.A(net572),
    .B(net502),
    .Y(_02087_));
 sky130_fd_sc_hd__nand2_1 _06787_ (.A(\core.CPU_Dmem_value_a5[4][24] ),
    .B(net447),
    .Y(_02088_));
 sky130_fd_sc_hd__a21oi_1 _06788_ (.A1(_02087_),
    .A2(_02088_),
    .B1(net601),
    .Y(_00544_));
 sky130_fd_sc_hd__nand2_1 _06789_ (.A(net571),
    .B(net502),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_1 _06790_ (.A(\core.CPU_Dmem_value_a5[4][25] ),
    .B(_02050_),
    .Y(_02090_));
 sky130_fd_sc_hd__a21oi_1 _06791_ (.A1(_02089_),
    .A2(_02090_),
    .B1(net601),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _06792_ (.A(net570),
    .B(net501),
    .Y(_02091_));
 sky130_fd_sc_hd__nand2_1 _06793_ (.A(\core.CPU_Dmem_value_a5[4][26] ),
    .B(net447),
    .Y(_02092_));
 sky130_fd_sc_hd__a21oi_1 _06794_ (.A1(_02091_),
    .A2(_02092_),
    .B1(net603),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _06796_ (.A(net569),
    .B(net501),
    .Y(_02094_));
 sky130_fd_sc_hd__nand2_1 _06798_ (.A(\core.CPU_Dmem_value_a5[4][27] ),
    .B(net447),
    .Y(_02096_));
 sky130_fd_sc_hd__a21oi_1 _06799_ (.A1(_02094_),
    .A2(_02096_),
    .B1(net604),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_1 _06800_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net502),
    .Y(_02097_));
 sky130_fd_sc_hd__nand2_1 _06801_ (.A(\core.CPU_Dmem_value_a5[4][28] ),
    .B(_02050_),
    .Y(_02098_));
 sky130_fd_sc_hd__a21oi_1 _06802_ (.A1(_02097_),
    .A2(_02098_),
    .B1(net600),
    .Y(_00548_));
 sky130_fd_sc_hd__nand2_1 _06803_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net502),
    .Y(_02099_));
 sky130_fd_sc_hd__nand2_1 _06804_ (.A(\core.CPU_Dmem_value_a5[4][29] ),
    .B(_02050_),
    .Y(_02100_));
 sky130_fd_sc_hd__a21oi_1 _06806_ (.A1(_02099_),
    .A2(_02100_),
    .B1(net602),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _06807_ (.A(\core.CPU_Dmem_value_a5[4][2] ),
    .B(net447),
    .Y(_02102_));
 sky130_fd_sc_hd__nand2_1 _06808_ (.A(net568),
    .B(net501),
    .Y(_02103_));
 sky130_fd_sc_hd__nand3b_1 _06809_ (.A_N(net605),
    .B(_02102_),
    .C(_02103_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _06810_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net502),
    .Y(_02104_));
 sky130_fd_sc_hd__nand2_1 _06811_ (.A(\core.CPU_Dmem_value_a5[4][30] ),
    .B(_02050_),
    .Y(_02105_));
 sky130_fd_sc_hd__a21oi_1 _06812_ (.A1(_02104_),
    .A2(_02105_),
    .B1(net602),
    .Y(_00551_));
 sky130_fd_sc_hd__nand2_1 _06813_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net501),
    .Y(_02106_));
 sky130_fd_sc_hd__nand2_1 _06814_ (.A(\core.CPU_Dmem_value_a5[4][31] ),
    .B(net447),
    .Y(_02107_));
 sky130_fd_sc_hd__a21oi_1 _06815_ (.A1(_02106_),
    .A2(_02107_),
    .B1(net601),
    .Y(_00552_));
 sky130_fd_sc_hd__nand2_1 _06816_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net502),
    .Y(_02108_));
 sky130_fd_sc_hd__nand2_1 _06817_ (.A(\core.CPU_Dmem_value_a5[4][3] ),
    .B(_02050_),
    .Y(_02109_));
 sky130_fd_sc_hd__a21oi_1 _06818_ (.A1(_02108_),
    .A2(_02109_),
    .B1(net602),
    .Y(_00553_));
 sky130_fd_sc_hd__nand2_1 _06819_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net501),
    .Y(_02110_));
 sky130_fd_sc_hd__nand2_1 _06820_ (.A(\core.CPU_Dmem_value_a5[4][4] ),
    .B(_02050_),
    .Y(_02111_));
 sky130_fd_sc_hd__a21oi_1 _06821_ (.A1(_02110_),
    .A2(_02111_),
    .B1(net599),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_1 _06822_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net501),
    .Y(_02112_));
 sky130_fd_sc_hd__nand2_1 _06823_ (.A(\core.CPU_Dmem_value_a5[4][5] ),
    .B(_02050_),
    .Y(_02113_));
 sky130_fd_sc_hd__a21oi_1 _06824_ (.A1(_02112_),
    .A2(_02113_),
    .B1(net605),
    .Y(_00555_));
 sky130_fd_sc_hd__nand2_1 _06825_ (.A(net567),
    .B(net502),
    .Y(_02114_));
 sky130_fd_sc_hd__nand2_1 _06826_ (.A(\core.CPU_Dmem_value_a5[4][6] ),
    .B(_02050_),
    .Y(_02115_));
 sky130_fd_sc_hd__a21oi_1 _06827_ (.A1(_02114_),
    .A2(_02115_),
    .B1(net599),
    .Y(_00556_));
 sky130_fd_sc_hd__nand2_1 _06828_ (.A(net566),
    .B(net502),
    .Y(_02116_));
 sky130_fd_sc_hd__nand2_1 _06829_ (.A(\core.CPU_Dmem_value_a5[4][7] ),
    .B(_02050_),
    .Y(_02117_));
 sky130_fd_sc_hd__a21oi_1 _06830_ (.A1(_02116_),
    .A2(_02117_),
    .B1(net599),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _06831_ (.A(net565),
    .B(net501),
    .Y(_02118_));
 sky130_fd_sc_hd__nand2_1 _06832_ (.A(\core.CPU_Dmem_value_a5[4][8] ),
    .B(net447),
    .Y(_02119_));
 sky130_fd_sc_hd__a21oi_1 _06833_ (.A1(_02118_),
    .A2(_02119_),
    .B1(net601),
    .Y(_00558_));
 sky130_fd_sc_hd__nand2_1 _06834_ (.A(net564),
    .B(net501),
    .Y(_02120_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(\core.CPU_Dmem_value_a5[4][9] ),
    .B(net447),
    .Y(_02121_));
 sky130_fd_sc_hd__a21oi_1 _06836_ (.A1(_02120_),
    .A2(_02121_),
    .B1(net603),
    .Y(_00559_));
 sky130_fd_sc_hd__nor2_4 _06837_ (.A(_01580_),
    .B(_02044_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_2 _06838_ (.A(net560),
    .B(net498),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(\core.CPU_Dmem_value_a5[5][0] ),
    .B(_02123_),
    .Y(_02125_));
 sky130_fd_sc_hd__nor3_2 _06841_ (.A(net561),
    .B(_01580_),
    .C(_02044_),
    .Y(_02126_));
 sky130_fd_sc_hd__nand2_1 _06843_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net496),
    .Y(_02128_));
 sky130_fd_sc_hd__nand3b_1 _06844_ (.A_N(\core.CPU_reset_a4 ),
    .B(_02125_),
    .C(_02128_),
    .Y(_00560_));
 sky130_fd_sc_hd__nand2_1 _06845_ (.A(net584),
    .B(net496),
    .Y(_02129_));
 sky130_fd_sc_hd__nand2_1 _06846_ (.A(\core.CPU_Dmem_value_a5[5][10] ),
    .B(net446),
    .Y(_02130_));
 sky130_fd_sc_hd__a21oi_1 _06848_ (.A1(_02129_),
    .A2(_02130_),
    .B1(net601),
    .Y(_00561_));
 sky130_fd_sc_hd__nand2_1 _06849_ (.A(net583),
    .B(net495),
    .Y(_02132_));
 sky130_fd_sc_hd__nand2_1 _06850_ (.A(\core.CPU_Dmem_value_a5[5][11] ),
    .B(net446),
    .Y(_02133_));
 sky130_fd_sc_hd__a21oi_1 _06851_ (.A1(_02132_),
    .A2(_02133_),
    .B1(net600),
    .Y(_00562_));
 sky130_fd_sc_hd__nand2_1 _06852_ (.A(net582),
    .B(net495),
    .Y(_02134_));
 sky130_fd_sc_hd__nand2_1 _06853_ (.A(\core.CPU_Dmem_value_a5[5][12] ),
    .B(net446),
    .Y(_02135_));
 sky130_fd_sc_hd__a21oi_1 _06854_ (.A1(_02134_),
    .A2(_02135_),
    .B1(net602),
    .Y(_00563_));
 sky130_fd_sc_hd__nand2_1 _06855_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net496),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_1 _06856_ (.A(\core.CPU_Dmem_value_a5[5][13] ),
    .B(net446),
    .Y(_02137_));
 sky130_fd_sc_hd__a21oi_1 _06857_ (.A1(_02136_),
    .A2(_02137_),
    .B1(net605),
    .Y(_00564_));
 sky130_fd_sc_hd__nand2_1 _06858_ (.A(net581),
    .B(net495),
    .Y(_02138_));
 sky130_fd_sc_hd__nand2_1 _06859_ (.A(\core.CPU_Dmem_value_a5[5][14] ),
    .B(net446),
    .Y(_02139_));
 sky130_fd_sc_hd__a21oi_1 _06860_ (.A1(_02138_),
    .A2(_02139_),
    .B1(net599),
    .Y(_00565_));
 sky130_fd_sc_hd__nand2_1 _06861_ (.A(net580),
    .B(net496),
    .Y(_02140_));
 sky130_fd_sc_hd__nand2_1 _06862_ (.A(\core.CPU_Dmem_value_a5[5][15] ),
    .B(net446),
    .Y(_02141_));
 sky130_fd_sc_hd__a21oi_1 _06863_ (.A1(_02140_),
    .A2(_02141_),
    .B1(net603),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _06864_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net496),
    .Y(_02142_));
 sky130_fd_sc_hd__nand2_1 _06865_ (.A(\core.CPU_Dmem_value_a5[5][16] ),
    .B(_02123_),
    .Y(_02143_));
 sky130_fd_sc_hd__a21oi_1 _06866_ (.A1(_02142_),
    .A2(_02143_),
    .B1(net604),
    .Y(_00567_));
 sky130_fd_sc_hd__nand2_1 _06867_ (.A(net579),
    .B(net496),
    .Y(_02144_));
 sky130_fd_sc_hd__nand2_1 _06868_ (.A(\core.CPU_Dmem_value_a5[5][17] ),
    .B(_02123_),
    .Y(_02145_));
 sky130_fd_sc_hd__a21oi_1 _06869_ (.A1(_02144_),
    .A2(_02145_),
    .B1(net604),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _06871_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net496),
    .Y(_02147_));
 sky130_fd_sc_hd__nand2_1 _06873_ (.A(\core.CPU_Dmem_value_a5[5][18] ),
    .B(_02123_),
    .Y(_02149_));
 sky130_fd_sc_hd__a21oi_1 _06874_ (.A1(_02147_),
    .A2(_02149_),
    .B1(net604),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _06875_ (.A(net578),
    .B(net495),
    .Y(_02150_));
 sky130_fd_sc_hd__nand2_1 _06876_ (.A(\core.CPU_Dmem_value_a5[5][19] ),
    .B(net446),
    .Y(_02151_));
 sky130_fd_sc_hd__a21oi_1 _06877_ (.A1(_02150_),
    .A2(_02151_),
    .B1(net600),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _06878_ (.A(net577),
    .B(net496),
    .Y(_02152_));
 sky130_fd_sc_hd__nand2_1 _06879_ (.A(\core.CPU_Dmem_value_a5[5][1] ),
    .B(net446),
    .Y(_02153_));
 sky130_fd_sc_hd__a21oi_1 _06881_ (.A1(_02152_),
    .A2(_02153_),
    .B1(net605),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _06882_ (.A(net576),
    .B(net495),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_1 _06883_ (.A(\core.CPU_Dmem_value_a5[5][20] ),
    .B(net446),
    .Y(_02156_));
 sky130_fd_sc_hd__a21oi_1 _06884_ (.A1(_02155_),
    .A2(_02156_),
    .B1(net601),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_1 _06885_ (.A(net575),
    .B(net496),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2_1 _06886_ (.A(\core.CPU_Dmem_value_a5[5][21] ),
    .B(net446),
    .Y(_02158_));
 sky130_fd_sc_hd__a21oi_1 _06887_ (.A1(_02157_),
    .A2(_02158_),
    .B1(net601),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _06888_ (.A(net574),
    .B(net495),
    .Y(_02159_));
 sky130_fd_sc_hd__nand2_1 _06889_ (.A(\core.CPU_Dmem_value_a5[5][22] ),
    .B(net446),
    .Y(_02160_));
 sky130_fd_sc_hd__a21oi_1 _06890_ (.A1(_02159_),
    .A2(_02160_),
    .B1(net601),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _06891_ (.A(net573),
    .B(net495),
    .Y(_02161_));
 sky130_fd_sc_hd__nand2_1 _06892_ (.A(\core.CPU_Dmem_value_a5[5][23] ),
    .B(net446),
    .Y(_02162_));
 sky130_fd_sc_hd__a21oi_1 _06893_ (.A1(_02161_),
    .A2(_02162_),
    .B1(net601),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _06894_ (.A(net572),
    .B(net495),
    .Y(_02163_));
 sky130_fd_sc_hd__nand2_1 _06895_ (.A(\core.CPU_Dmem_value_a5[5][24] ),
    .B(net446),
    .Y(_02164_));
 sky130_fd_sc_hd__a21oi_1 _06896_ (.A1(_02163_),
    .A2(_02164_),
    .B1(net600),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2_1 _06897_ (.A(net571),
    .B(net495),
    .Y(_02165_));
 sky130_fd_sc_hd__nand2_1 _06898_ (.A(\core.CPU_Dmem_value_a5[5][25] ),
    .B(net446),
    .Y(_02166_));
 sky130_fd_sc_hd__a21oi_1 _06899_ (.A1(_02165_),
    .A2(_02166_),
    .B1(net601),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _06900_ (.A(net570),
    .B(net496),
    .Y(_02167_));
 sky130_fd_sc_hd__nand2_1 _06901_ (.A(\core.CPU_Dmem_value_a5[5][26] ),
    .B(net446),
    .Y(_02168_));
 sky130_fd_sc_hd__a21oi_1 _06902_ (.A1(_02167_),
    .A2(_02168_),
    .B1(net603),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _06904_ (.A(net569),
    .B(net496),
    .Y(_02170_));
 sky130_fd_sc_hd__nand2_1 _06906_ (.A(\core.CPU_Dmem_value_a5[5][27] ),
    .B(_02123_),
    .Y(_02172_));
 sky130_fd_sc_hd__a21oi_1 _06907_ (.A1(_02170_),
    .A2(_02172_),
    .B1(net604),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _06908_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net496),
    .Y(_02173_));
 sky130_fd_sc_hd__nand2_1 _06909_ (.A(\core.CPU_Dmem_value_a5[5][28] ),
    .B(_02123_),
    .Y(_02174_));
 sky130_fd_sc_hd__a21oi_1 _06910_ (.A1(_02173_),
    .A2(_02174_),
    .B1(net603),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2_1 _06911_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net495),
    .Y(_02175_));
 sky130_fd_sc_hd__nand2_1 _06912_ (.A(\core.CPU_Dmem_value_a5[5][29] ),
    .B(net446),
    .Y(_02176_));
 sky130_fd_sc_hd__a21oi_1 _06914_ (.A1(_02175_),
    .A2(_02176_),
    .B1(net599),
    .Y(_00581_));
 sky130_fd_sc_hd__nand2_1 _06915_ (.A(\core.CPU_Dmem_value_a5[5][2] ),
    .B(net446),
    .Y(_02178_));
 sky130_fd_sc_hd__nand2_1 _06916_ (.A(net568),
    .B(net496),
    .Y(_02179_));
 sky130_fd_sc_hd__nand3b_1 _06917_ (.A_N(net605),
    .B(_02178_),
    .C(_02179_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand2_1 _06918_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net495),
    .Y(_02180_));
 sky130_fd_sc_hd__nand2_1 _06919_ (.A(\core.CPU_Dmem_value_a5[5][30] ),
    .B(net446),
    .Y(_02181_));
 sky130_fd_sc_hd__a21oi_1 _06920_ (.A1(_02180_),
    .A2(_02181_),
    .B1(net599),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _06921_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net496),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_1 _06922_ (.A(\core.CPU_Dmem_value_a5[5][31] ),
    .B(net446),
    .Y(_02183_));
 sky130_fd_sc_hd__a21oi_1 _06923_ (.A1(_02182_),
    .A2(_02183_),
    .B1(net601),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _06924_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net496),
    .Y(_02184_));
 sky130_fd_sc_hd__nand2_1 _06925_ (.A(\core.CPU_Dmem_value_a5[5][3] ),
    .B(_02123_),
    .Y(_02185_));
 sky130_fd_sc_hd__a21oi_1 _06926_ (.A1(_02184_),
    .A2(_02185_),
    .B1(net600),
    .Y(_00585_));
 sky130_fd_sc_hd__nand2_1 _06927_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net496),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _06928_ (.A(\core.CPU_Dmem_value_a5[5][4] ),
    .B(_02123_),
    .Y(_02187_));
 sky130_fd_sc_hd__a21oi_1 _06929_ (.A1(_02186_),
    .A2(_02187_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _06930_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net496),
    .Y(_02188_));
 sky130_fd_sc_hd__nand2_1 _06931_ (.A(\core.CPU_Dmem_value_a5[5][5] ),
    .B(_02123_),
    .Y(_02189_));
 sky130_fd_sc_hd__a21oi_1 _06932_ (.A1(_02188_),
    .A2(_02189_),
    .B1(net605),
    .Y(_00587_));
 sky130_fd_sc_hd__nand2_1 _06933_ (.A(net567),
    .B(net495),
    .Y(_02190_));
 sky130_fd_sc_hd__nand2_1 _06934_ (.A(\core.CPU_Dmem_value_a5[5][6] ),
    .B(net446),
    .Y(_02191_));
 sky130_fd_sc_hd__a21oi_1 _06935_ (.A1(_02190_),
    .A2(_02191_),
    .B1(net599),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _06936_ (.A(net566),
    .B(net495),
    .Y(_02192_));
 sky130_fd_sc_hd__nand2_1 _06937_ (.A(\core.CPU_Dmem_value_a5[5][7] ),
    .B(net446),
    .Y(_02193_));
 sky130_fd_sc_hd__a21oi_1 _06938_ (.A1(_02192_),
    .A2(_02193_),
    .B1(net599),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_1 _06939_ (.A(net565),
    .B(net496),
    .Y(_02194_));
 sky130_fd_sc_hd__nand2_1 _06940_ (.A(\core.CPU_Dmem_value_a5[5][8] ),
    .B(net446),
    .Y(_02195_));
 sky130_fd_sc_hd__a21oi_1 _06941_ (.A1(_02194_),
    .A2(_02195_),
    .B1(net601),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _06942_ (.A(net564),
    .B(net496),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _06943_ (.A(\core.CPU_Dmem_value_a5[5][9] ),
    .B(net446),
    .Y(_02197_));
 sky130_fd_sc_hd__a21oi_1 _06944_ (.A1(_02196_),
    .A2(_02197_),
    .B1(net603),
    .Y(_00591_));
 sky130_fd_sc_hd__nor3_2 _06945_ (.A(net561),
    .B(_01344_),
    .C(_02044_),
    .Y(_02198_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net494),
    .Y(_02200_));
 sky130_fd_sc_hd__nor2_4 _06948_ (.A(_01344_),
    .B(_02044_),
    .Y(_02201_));
 sky130_fd_sc_hd__nand2_2 _06949_ (.A(net560),
    .B(net491),
    .Y(_02202_));
 sky130_fd_sc_hd__nand2_1 _06951_ (.A(\core.CPU_Dmem_value_a5[6][0] ),
    .B(_02202_),
    .Y(_02204_));
 sky130_fd_sc_hd__a21oi_1 _06953_ (.A1(_02200_),
    .A2(_02204_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00592_));
 sky130_fd_sc_hd__nand2_1 _06954_ (.A(net584),
    .B(net494),
    .Y(_02206_));
 sky130_fd_sc_hd__nand2_1 _06955_ (.A(\core.CPU_Dmem_value_a5[6][10] ),
    .B(net445),
    .Y(_02207_));
 sky130_fd_sc_hd__a21oi_1 _06956_ (.A1(_02206_),
    .A2(_02207_),
    .B1(net601),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _06957_ (.A(net583),
    .B(net493),
    .Y(_02208_));
 sky130_fd_sc_hd__nand2_1 _06958_ (.A(\core.CPU_Dmem_value_a5[6][11] ),
    .B(net445),
    .Y(_02209_));
 sky130_fd_sc_hd__a21oi_1 _06959_ (.A1(_02208_),
    .A2(_02209_),
    .B1(net600),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_1 _06960_ (.A(net582),
    .B(net493),
    .Y(_02210_));
 sky130_fd_sc_hd__nand2_1 _06961_ (.A(\core.CPU_Dmem_value_a5[6][12] ),
    .B(net445),
    .Y(_02211_));
 sky130_fd_sc_hd__a21oi_1 _06962_ (.A1(_02210_),
    .A2(_02211_),
    .B1(net602),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_1 _06963_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net494),
    .Y(_02212_));
 sky130_fd_sc_hd__nand2_1 _06964_ (.A(\core.CPU_Dmem_value_a5[6][13] ),
    .B(_02202_),
    .Y(_02213_));
 sky130_fd_sc_hd__a21oi_1 _06965_ (.A1(_02212_),
    .A2(_02213_),
    .B1(net605),
    .Y(_00596_));
 sky130_fd_sc_hd__nand2_1 _06966_ (.A(net581),
    .B(net493),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_1 _06967_ (.A(\core.CPU_Dmem_value_a5[6][14] ),
    .B(net445),
    .Y(_02215_));
 sky130_fd_sc_hd__a21oi_1 _06968_ (.A1(_02214_),
    .A2(_02215_),
    .B1(net599),
    .Y(_00597_));
 sky130_fd_sc_hd__nand2_1 _06969_ (.A(net580),
    .B(net494),
    .Y(_02216_));
 sky130_fd_sc_hd__nand2_1 _06970_ (.A(\core.CPU_Dmem_value_a5[6][15] ),
    .B(net445),
    .Y(_02217_));
 sky130_fd_sc_hd__a21oi_1 _06971_ (.A1(_02216_),
    .A2(_02217_),
    .B1(net601),
    .Y(_00598_));
 sky130_fd_sc_hd__nand2_1 _06972_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net494),
    .Y(_02218_));
 sky130_fd_sc_hd__nand2_1 _06973_ (.A(\core.CPU_Dmem_value_a5[6][16] ),
    .B(_02202_),
    .Y(_02219_));
 sky130_fd_sc_hd__a21oi_1 _06974_ (.A1(_02218_),
    .A2(_02219_),
    .B1(net603),
    .Y(_00599_));
 sky130_fd_sc_hd__nand2_1 _06976_ (.A(net579),
    .B(net494),
    .Y(_02221_));
 sky130_fd_sc_hd__nand2_1 _06978_ (.A(\core.CPU_Dmem_value_a5[6][17] ),
    .B(_02202_),
    .Y(_02223_));
 sky130_fd_sc_hd__a21oi_1 _06979_ (.A1(_02221_),
    .A2(_02223_),
    .B1(net604),
    .Y(_00600_));
 sky130_fd_sc_hd__nand2_1 _06980_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net494),
    .Y(_02224_));
 sky130_fd_sc_hd__nand2_1 _06981_ (.A(\core.CPU_Dmem_value_a5[6][18] ),
    .B(_02202_),
    .Y(_02225_));
 sky130_fd_sc_hd__a21oi_1 _06982_ (.A1(_02224_),
    .A2(_02225_),
    .B1(net604),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_1 _06983_ (.A(net578),
    .B(net493),
    .Y(_02226_));
 sky130_fd_sc_hd__nand2_1 _06984_ (.A(\core.CPU_Dmem_value_a5[6][19] ),
    .B(net445),
    .Y(_02227_));
 sky130_fd_sc_hd__a21oi_1 _06986_ (.A1(_02226_),
    .A2(_02227_),
    .B1(net600),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2_1 _06987_ (.A(\core.CPU_Dmem_value_a5[6][1] ),
    .B(_02202_),
    .Y(_02229_));
 sky130_fd_sc_hd__nand2_1 _06988_ (.A(net577),
    .B(net494),
    .Y(_02230_));
 sky130_fd_sc_hd__nand3b_1 _06989_ (.A_N(net605),
    .B(_02229_),
    .C(_02230_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _06990_ (.A(net576),
    .B(net494),
    .Y(_02231_));
 sky130_fd_sc_hd__nand2_1 _06991_ (.A(\core.CPU_Dmem_value_a5[6][20] ),
    .B(_02202_),
    .Y(_02232_));
 sky130_fd_sc_hd__a21oi_1 _06992_ (.A1(_02231_),
    .A2(_02232_),
    .B1(net601),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _06993_ (.A(net575),
    .B(net494),
    .Y(_02233_));
 sky130_fd_sc_hd__nand2_1 _06994_ (.A(\core.CPU_Dmem_value_a5[6][21] ),
    .B(_02202_),
    .Y(_02234_));
 sky130_fd_sc_hd__a21oi_1 _06995_ (.A1(_02233_),
    .A2(_02234_),
    .B1(net605),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_1 _06996_ (.A(net574),
    .B(net494),
    .Y(_02235_));
 sky130_fd_sc_hd__nand2_1 _06997_ (.A(\core.CPU_Dmem_value_a5[6][22] ),
    .B(net445),
    .Y(_02236_));
 sky130_fd_sc_hd__a21oi_1 _06998_ (.A1(_02235_),
    .A2(_02236_),
    .B1(net601),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_1 _06999_ (.A(net573),
    .B(net493),
    .Y(_02237_));
 sky130_fd_sc_hd__nand2_1 _07000_ (.A(\core.CPU_Dmem_value_a5[6][23] ),
    .B(net445),
    .Y(_02238_));
 sky130_fd_sc_hd__a21oi_1 _07001_ (.A1(_02237_),
    .A2(_02238_),
    .B1(net601),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_1 _07002_ (.A(net572),
    .B(net494),
    .Y(_02239_));
 sky130_fd_sc_hd__nand2_1 _07003_ (.A(\core.CPU_Dmem_value_a5[6][24] ),
    .B(net445),
    .Y(_02240_));
 sky130_fd_sc_hd__a21oi_1 _07004_ (.A1(_02239_),
    .A2(_02240_),
    .B1(net601),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _07005_ (.A(net571),
    .B(net494),
    .Y(_02241_));
 sky130_fd_sc_hd__nand2_1 _07006_ (.A(\core.CPU_Dmem_value_a5[6][25] ),
    .B(_02202_),
    .Y(_02242_));
 sky130_fd_sc_hd__a21oi_1 _07007_ (.A1(_02241_),
    .A2(_02242_),
    .B1(net601),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_1 _07008_ (.A(net570),
    .B(net494),
    .Y(_02243_));
 sky130_fd_sc_hd__nand2_1 _07009_ (.A(\core.CPU_Dmem_value_a5[6][26] ),
    .B(_02202_),
    .Y(_02244_));
 sky130_fd_sc_hd__a21oi_1 _07010_ (.A1(_02243_),
    .A2(_02244_),
    .B1(net603),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_1 _07012_ (.A(net569),
    .B(net494),
    .Y(_02246_));
 sky130_fd_sc_hd__nand2_1 _07014_ (.A(\core.CPU_Dmem_value_a5[6][27] ),
    .B(_02202_),
    .Y(_02248_));
 sky130_fd_sc_hd__a21oi_1 _07015_ (.A1(_02246_),
    .A2(_02248_),
    .B1(net604),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _07016_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net494),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_1 _07017_ (.A(\core.CPU_Dmem_value_a5[6][28] ),
    .B(_02202_),
    .Y(_02250_));
 sky130_fd_sc_hd__a21oi_1 _07018_ (.A1(_02249_),
    .A2(_02250_),
    .B1(net603),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _07019_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net493),
    .Y(_02251_));
 sky130_fd_sc_hd__nand2_1 _07020_ (.A(\core.CPU_Dmem_value_a5[6][29] ),
    .B(net445),
    .Y(_02252_));
 sky130_fd_sc_hd__a21oi_1 _07023_ (.A1(_02251_),
    .A2(_02252_),
    .B1(net599),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _07024_ (.A(\core.CPU_Dmem_value_a5[6][2] ),
    .B(_02202_),
    .Y(_02255_));
 sky130_fd_sc_hd__nand2_1 _07025_ (.A(net568),
    .B(net494),
    .Y(_02256_));
 sky130_fd_sc_hd__nand3b_1 _07026_ (.A_N(net605),
    .B(_02255_),
    .C(_02256_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_1 _07027_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net493),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_1 _07028_ (.A(\core.CPU_Dmem_value_a5[6][30] ),
    .B(net445),
    .Y(_02258_));
 sky130_fd_sc_hd__a21oi_1 _07029_ (.A1(_02257_),
    .A2(_02258_),
    .B1(net599),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2_1 _07030_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net494),
    .Y(_02259_));
 sky130_fd_sc_hd__nand2_1 _07031_ (.A(\core.CPU_Dmem_value_a5[6][31] ),
    .B(net445),
    .Y(_02260_));
 sky130_fd_sc_hd__a21oi_1 _07032_ (.A1(_02259_),
    .A2(_02260_),
    .B1(net601),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_1 _07033_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net493),
    .Y(_02261_));
 sky130_fd_sc_hd__nand2_1 _07034_ (.A(\core.CPU_Dmem_value_a5[6][3] ),
    .B(net445),
    .Y(_02262_));
 sky130_fd_sc_hd__a21oi_1 _07035_ (.A1(_02261_),
    .A2(_02262_),
    .B1(net599),
    .Y(_00617_));
 sky130_fd_sc_hd__nand2_1 _07036_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net493),
    .Y(_02263_));
 sky130_fd_sc_hd__nand2_1 _07037_ (.A(\core.CPU_Dmem_value_a5[6][4] ),
    .B(_02202_),
    .Y(_02264_));
 sky130_fd_sc_hd__a21oi_1 _07038_ (.A1(_02263_),
    .A2(_02264_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00618_));
 sky130_fd_sc_hd__nand2_1 _07039_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net494),
    .Y(_02265_));
 sky130_fd_sc_hd__nand2_1 _07040_ (.A(\core.CPU_Dmem_value_a5[6][5] ),
    .B(_02202_),
    .Y(_02266_));
 sky130_fd_sc_hd__a21oi_1 _07041_ (.A1(_02265_),
    .A2(_02266_),
    .B1(net605),
    .Y(_00619_));
 sky130_fd_sc_hd__nand2_1 _07042_ (.A(net567),
    .B(net493),
    .Y(_02267_));
 sky130_fd_sc_hd__nand2_1 _07043_ (.A(\core.CPU_Dmem_value_a5[6][6] ),
    .B(net445),
    .Y(_02268_));
 sky130_fd_sc_hd__a21oi_1 _07044_ (.A1(_02267_),
    .A2(_02268_),
    .B1(net599),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2_1 _07045_ (.A(net566),
    .B(net493),
    .Y(_02269_));
 sky130_fd_sc_hd__nand2_1 _07046_ (.A(\core.CPU_Dmem_value_a5[6][7] ),
    .B(net445),
    .Y(_02270_));
 sky130_fd_sc_hd__a21oi_1 _07047_ (.A1(_02269_),
    .A2(_02270_),
    .B1(net602),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _07048_ (.A(net565),
    .B(net494),
    .Y(_02271_));
 sky130_fd_sc_hd__nand2_1 _07049_ (.A(\core.CPU_Dmem_value_a5[6][8] ),
    .B(net445),
    .Y(_02272_));
 sky130_fd_sc_hd__a21oi_1 _07050_ (.A1(_02271_),
    .A2(_02272_),
    .B1(net601),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _07051_ (.A(net564),
    .B(net494),
    .Y(_02273_));
 sky130_fd_sc_hd__nand2_1 _07052_ (.A(\core.CPU_Dmem_value_a5[6][9] ),
    .B(_02202_),
    .Y(_02274_));
 sky130_fd_sc_hd__a21oi_1 _07053_ (.A1(_02273_),
    .A2(_02274_),
    .B1(net605),
    .Y(_00623_));
 sky130_fd_sc_hd__nor2_4 _07054_ (.A(_01425_),
    .B(_02044_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand2_2 _07056_ (.A(net560),
    .B(_02275_),
    .Y(_02277_));
 sky130_fd_sc_hd__nand2_1 _07058_ (.A(\core.CPU_Dmem_value_a5[7][0] ),
    .B(net444),
    .Y(_02279_));
 sky130_fd_sc_hd__nor3_2 _07059_ (.A(net561),
    .B(_01425_),
    .C(_02044_),
    .Y(_02280_));
 sky130_fd_sc_hd__nand2_1 _07061_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net489),
    .Y(_02282_));
 sky130_fd_sc_hd__nand3b_1 _07062_ (.A_N(\core.CPU_reset_a4 ),
    .B(_02279_),
    .C(_02282_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _07063_ (.A(net584),
    .B(net489),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _07064_ (.A(\core.CPU_Dmem_value_a5[7][10] ),
    .B(_02277_),
    .Y(_02284_));
 sky130_fd_sc_hd__a21oi_1 _07066_ (.A1(_02283_),
    .A2(_02284_),
    .B1(net601),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _07067_ (.A(net583),
    .B(net489),
    .Y(_02286_));
 sky130_fd_sc_hd__nand2_1 _07068_ (.A(\core.CPU_Dmem_value_a5[7][11] ),
    .B(net444),
    .Y(_02287_));
 sky130_fd_sc_hd__a21oi_1 _07069_ (.A1(_02286_),
    .A2(_02287_),
    .B1(net600),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _07070_ (.A(net582),
    .B(net488),
    .Y(_02288_));
 sky130_fd_sc_hd__nand2_1 _07071_ (.A(\core.CPU_Dmem_value_a5[7][12] ),
    .B(net444),
    .Y(_02289_));
 sky130_fd_sc_hd__a21oi_1 _07072_ (.A1(_02288_),
    .A2(_02289_),
    .B1(net602),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _07073_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net489),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_1 _07074_ (.A(\core.CPU_Dmem_value_a5[7][13] ),
    .B(_02277_),
    .Y(_02291_));
 sky130_fd_sc_hd__a21oi_1 _07075_ (.A1(_02290_),
    .A2(_02291_),
    .B1(net604),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _07076_ (.A(net581),
    .B(net488),
    .Y(_02292_));
 sky130_fd_sc_hd__nand2_1 _07077_ (.A(\core.CPU_Dmem_value_a5[7][14] ),
    .B(net444),
    .Y(_02293_));
 sky130_fd_sc_hd__a21oi_1 _07078_ (.A1(_02292_),
    .A2(_02293_),
    .B1(net599),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_1 _07079_ (.A(net580),
    .B(net489),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_1 _07080_ (.A(\core.CPU_Dmem_value_a5[7][15] ),
    .B(_02277_),
    .Y(_02295_));
 sky130_fd_sc_hd__a21oi_1 _07081_ (.A1(_02294_),
    .A2(_02295_),
    .B1(net603),
    .Y(_00630_));
 sky130_fd_sc_hd__nand2_1 _07082_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net489),
    .Y(_02296_));
 sky130_fd_sc_hd__nand2_1 _07083_ (.A(\core.CPU_Dmem_value_a5[7][16] ),
    .B(net444),
    .Y(_02297_));
 sky130_fd_sc_hd__a21oi_1 _07084_ (.A1(_02296_),
    .A2(_02297_),
    .B1(net603),
    .Y(_00631_));
 sky130_fd_sc_hd__nand2_1 _07086_ (.A(net579),
    .B(net489),
    .Y(_02299_));
 sky130_fd_sc_hd__nand2_1 _07088_ (.A(\core.CPU_Dmem_value_a5[7][17] ),
    .B(_02277_),
    .Y(_02301_));
 sky130_fd_sc_hd__a21oi_1 _07089_ (.A1(_02299_),
    .A2(_02301_),
    .B1(net604),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _07090_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net489),
    .Y(_02302_));
 sky130_fd_sc_hd__nand2_1 _07091_ (.A(\core.CPU_Dmem_value_a5[7][18] ),
    .B(net444),
    .Y(_02303_));
 sky130_fd_sc_hd__a21oi_1 _07092_ (.A1(_02302_),
    .A2(_02303_),
    .B1(net604),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _07093_ (.A(net578),
    .B(net489),
    .Y(_02304_));
 sky130_fd_sc_hd__nand2_1 _07094_ (.A(\core.CPU_Dmem_value_a5[7][19] ),
    .B(net444),
    .Y(_02305_));
 sky130_fd_sc_hd__a21oi_1 _07095_ (.A1(_02304_),
    .A2(_02305_),
    .B1(net600),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _07096_ (.A(\core.CPU_Dmem_value_a5[7][1] ),
    .B(_02277_),
    .Y(_02306_));
 sky130_fd_sc_hd__nand2_1 _07097_ (.A(net577),
    .B(net489),
    .Y(_02307_));
 sky130_fd_sc_hd__nand3b_1 _07098_ (.A_N(net605),
    .B(_02306_),
    .C(_02307_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _07099_ (.A(net576),
    .B(net489),
    .Y(_02308_));
 sky130_fd_sc_hd__nand2_1 _07100_ (.A(\core.CPU_Dmem_value_a5[7][20] ),
    .B(_02277_),
    .Y(_02309_));
 sky130_fd_sc_hd__a21oi_1 _07102_ (.A1(_02308_),
    .A2(_02309_),
    .B1(net601),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _07103_ (.A(net575),
    .B(net489),
    .Y(_02311_));
 sky130_fd_sc_hd__nand2_1 _07104_ (.A(\core.CPU_Dmem_value_a5[7][21] ),
    .B(_02277_),
    .Y(_02312_));
 sky130_fd_sc_hd__a21oi_1 _07105_ (.A1(_02311_),
    .A2(_02312_),
    .B1(net603),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_1 _07106_ (.A(net574),
    .B(net489),
    .Y(_02313_));
 sky130_fd_sc_hd__nand2_1 _07107_ (.A(\core.CPU_Dmem_value_a5[7][22] ),
    .B(_02277_),
    .Y(_02314_));
 sky130_fd_sc_hd__a21oi_1 _07108_ (.A1(_02313_),
    .A2(_02314_),
    .B1(net601),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _07109_ (.A(net573),
    .B(net489),
    .Y(_02315_));
 sky130_fd_sc_hd__nand2_1 _07110_ (.A(\core.CPU_Dmem_value_a5[7][23] ),
    .B(_02277_),
    .Y(_02316_));
 sky130_fd_sc_hd__a21oi_1 _07111_ (.A1(_02315_),
    .A2(_02316_),
    .B1(net601),
    .Y(_00639_));
 sky130_fd_sc_hd__nand2_1 _07112_ (.A(net572),
    .B(net489),
    .Y(_02317_));
 sky130_fd_sc_hd__nand2_1 _07113_ (.A(\core.CPU_Dmem_value_a5[7][24] ),
    .B(net444),
    .Y(_02318_));
 sky130_fd_sc_hd__a21oi_1 _07114_ (.A1(_02317_),
    .A2(_02318_),
    .B1(net600),
    .Y(_00640_));
 sky130_fd_sc_hd__nand2_1 _07115_ (.A(net571),
    .B(net489),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_1 _07116_ (.A(\core.CPU_Dmem_value_a5[7][25] ),
    .B(net444),
    .Y(_02320_));
 sky130_fd_sc_hd__a21oi_1 _07117_ (.A1(_02319_),
    .A2(_02320_),
    .B1(net601),
    .Y(_00641_));
 sky130_fd_sc_hd__nand2_1 _07118_ (.A(net570),
    .B(net489),
    .Y(_02321_));
 sky130_fd_sc_hd__nand2_1 _07119_ (.A(\core.CPU_Dmem_value_a5[7][26] ),
    .B(_02277_),
    .Y(_02322_));
 sky130_fd_sc_hd__a21oi_1 _07120_ (.A1(_02321_),
    .A2(_02322_),
    .B1(net603),
    .Y(_00642_));
 sky130_fd_sc_hd__nand2_1 _07122_ (.A(net569),
    .B(net489),
    .Y(_02324_));
 sky130_fd_sc_hd__nand2_1 _07124_ (.A(\core.CPU_Dmem_value_a5[7][27] ),
    .B(_02277_),
    .Y(_02326_));
 sky130_fd_sc_hd__a21oi_1 _07125_ (.A1(_02324_),
    .A2(_02326_),
    .B1(net604),
    .Y(_00643_));
 sky130_fd_sc_hd__nand2_1 _07126_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net489),
    .Y(_02327_));
 sky130_fd_sc_hd__nand2_1 _07127_ (.A(\core.CPU_Dmem_value_a5[7][28] ),
    .B(net444),
    .Y(_02328_));
 sky130_fd_sc_hd__a21oi_1 _07128_ (.A1(_02327_),
    .A2(_02328_),
    .B1(net600),
    .Y(_00644_));
 sky130_fd_sc_hd__nand2_1 _07129_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net488),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _07130_ (.A(\core.CPU_Dmem_value_a5[7][29] ),
    .B(net444),
    .Y(_02330_));
 sky130_fd_sc_hd__a21oi_1 _07131_ (.A1(_02329_),
    .A2(_02330_),
    .B1(net599),
    .Y(_00645_));
 sky130_fd_sc_hd__nand2_1 _07132_ (.A(\core.CPU_Dmem_value_a5[7][2] ),
    .B(_02277_),
    .Y(_02331_));
 sky130_fd_sc_hd__nand2_1 _07133_ (.A(net568),
    .B(net489),
    .Y(_02332_));
 sky130_fd_sc_hd__nand3b_1 _07134_ (.A_N(net605),
    .B(_02331_),
    .C(_02332_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand2_1 _07135_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net488),
    .Y(_02333_));
 sky130_fd_sc_hd__nand2_1 _07136_ (.A(\core.CPU_Dmem_value_a5[7][30] ),
    .B(net444),
    .Y(_02334_));
 sky130_fd_sc_hd__a21oi_1 _07138_ (.A1(_02333_),
    .A2(_02334_),
    .B1(net602),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2_1 _07139_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net489),
    .Y(_02336_));
 sky130_fd_sc_hd__nand2_1 _07140_ (.A(\core.CPU_Dmem_value_a5[7][31] ),
    .B(_02277_),
    .Y(_02337_));
 sky130_fd_sc_hd__a21oi_1 _07141_ (.A1(_02336_),
    .A2(_02337_),
    .B1(net601),
    .Y(_00648_));
 sky130_fd_sc_hd__nand2_1 _07142_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net489),
    .Y(_02338_));
 sky130_fd_sc_hd__nand2_1 _07143_ (.A(\core.CPU_Dmem_value_a5[7][3] ),
    .B(net444),
    .Y(_02339_));
 sky130_fd_sc_hd__a21oi_1 _07144_ (.A1(_02338_),
    .A2(_02339_),
    .B1(net600),
    .Y(_00649_));
 sky130_fd_sc_hd__nand2_1 _07145_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net489),
    .Y(_02340_));
 sky130_fd_sc_hd__nand2_1 _07146_ (.A(\core.CPU_Dmem_value_a5[7][4] ),
    .B(net444),
    .Y(_02341_));
 sky130_fd_sc_hd__a21oi_1 _07147_ (.A1(_02340_),
    .A2(_02341_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00650_));
 sky130_fd_sc_hd__nand2_1 _07148_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net489),
    .Y(_02342_));
 sky130_fd_sc_hd__nand2_1 _07149_ (.A(\core.CPU_Dmem_value_a5[7][5] ),
    .B(_02277_),
    .Y(_02343_));
 sky130_fd_sc_hd__a21oi_1 _07150_ (.A1(_02342_),
    .A2(_02343_),
    .B1(net605),
    .Y(_00651_));
 sky130_fd_sc_hd__nand2_1 _07151_ (.A(net567),
    .B(net488),
    .Y(_02344_));
 sky130_fd_sc_hd__nand2_1 _07152_ (.A(\core.CPU_Dmem_value_a5[7][6] ),
    .B(net444),
    .Y(_02345_));
 sky130_fd_sc_hd__a21oi_1 _07153_ (.A1(_02344_),
    .A2(_02345_),
    .B1(net599),
    .Y(_00652_));
 sky130_fd_sc_hd__nand2_1 _07154_ (.A(net566),
    .B(net488),
    .Y(_02346_));
 sky130_fd_sc_hd__nand2_1 _07155_ (.A(\core.CPU_Dmem_value_a5[7][7] ),
    .B(net444),
    .Y(_02347_));
 sky130_fd_sc_hd__a21oi_1 _07156_ (.A1(_02346_),
    .A2(_02347_),
    .B1(net599),
    .Y(_00653_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(net565),
    .B(net489),
    .Y(_02348_));
 sky130_fd_sc_hd__nand2_1 _07158_ (.A(\core.CPU_Dmem_value_a5[7][8] ),
    .B(_02277_),
    .Y(_02349_));
 sky130_fd_sc_hd__a21oi_1 _07159_ (.A1(_02348_),
    .A2(_02349_),
    .B1(net601),
    .Y(_00654_));
 sky130_fd_sc_hd__nand2_1 _07160_ (.A(net564),
    .B(net489),
    .Y(_02350_));
 sky130_fd_sc_hd__nand2_1 _07161_ (.A(\core.CPU_Dmem_value_a5[7][9] ),
    .B(_02277_),
    .Y(_02351_));
 sky130_fd_sc_hd__a21oi_1 _07162_ (.A1(_02350_),
    .A2(_02351_),
    .B1(net603),
    .Y(_00655_));
 sky130_fd_sc_hd__nor4_2 _07163_ (.A(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .C(net561),
    .D(_01346_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand2_1 _07165_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net486),
    .Y(_02354_));
 sky130_fd_sc_hd__nor3_2 _07166_ (.A(\core.CPU_dmem_addr_a4[1] ),
    .B(\core.CPU_dmem_addr_a4[0] ),
    .C(_01346_),
    .Y(_02355_));
 sky130_fd_sc_hd__nand2_2 _07167_ (.A(net560),
    .B(net485),
    .Y(_02356_));
 sky130_fd_sc_hd__nand2_1 _07169_ (.A(\core.CPU_Dmem_value_a5[8][0] ),
    .B(_02356_),
    .Y(_02358_));
 sky130_fd_sc_hd__a21oi_1 _07170_ (.A1(_02354_),
    .A2(_02358_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00656_));
 sky130_fd_sc_hd__nand2_1 _07171_ (.A(net584),
    .B(net487),
    .Y(_02359_));
 sky130_fd_sc_hd__nand2_1 _07172_ (.A(\core.CPU_Dmem_value_a5[8][10] ),
    .B(net443),
    .Y(_02360_));
 sky130_fd_sc_hd__a21oi_1 _07174_ (.A1(_02359_),
    .A2(_02360_),
    .B1(net601),
    .Y(_00657_));
 sky130_fd_sc_hd__nand2_1 _07175_ (.A(net583),
    .B(net487),
    .Y(_02362_));
 sky130_fd_sc_hd__nand2_1 _07176_ (.A(\core.CPU_Dmem_value_a5[8][11] ),
    .B(net443),
    .Y(_02363_));
 sky130_fd_sc_hd__a21oi_1 _07177_ (.A1(_02362_),
    .A2(_02363_),
    .B1(net600),
    .Y(_00658_));
 sky130_fd_sc_hd__nand2_1 _07178_ (.A(net582),
    .B(net487),
    .Y(_02364_));
 sky130_fd_sc_hd__nand2_1 _07179_ (.A(\core.CPU_Dmem_value_a5[8][12] ),
    .B(net443),
    .Y(_02365_));
 sky130_fd_sc_hd__a21oi_1 _07180_ (.A1(_02364_),
    .A2(_02365_),
    .B1(net600),
    .Y(_00659_));
 sky130_fd_sc_hd__nand2_1 _07181_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net486),
    .Y(_02366_));
 sky130_fd_sc_hd__nand2_1 _07182_ (.A(\core.CPU_Dmem_value_a5[8][13] ),
    .B(net443),
    .Y(_02367_));
 sky130_fd_sc_hd__a21oi_1 _07183_ (.A1(_02366_),
    .A2(_02367_),
    .B1(net604),
    .Y(_00660_));
 sky130_fd_sc_hd__nand2_1 _07184_ (.A(net581),
    .B(net487),
    .Y(_02368_));
 sky130_fd_sc_hd__nand2_1 _07185_ (.A(\core.CPU_Dmem_value_a5[8][14] ),
    .B(_02356_),
    .Y(_02369_));
 sky130_fd_sc_hd__a21oi_1 _07186_ (.A1(_02368_),
    .A2(_02369_),
    .B1(net599),
    .Y(_00661_));
 sky130_fd_sc_hd__nand2_1 _07187_ (.A(net580),
    .B(net487),
    .Y(_02370_));
 sky130_fd_sc_hd__nand2_1 _07188_ (.A(\core.CPU_Dmem_value_a5[8][15] ),
    .B(net443),
    .Y(_02371_));
 sky130_fd_sc_hd__a21oi_1 _07189_ (.A1(_02370_),
    .A2(_02371_),
    .B1(net601),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _07190_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net486),
    .Y(_02372_));
 sky130_fd_sc_hd__nand2_1 _07191_ (.A(\core.CPU_Dmem_value_a5[8][16] ),
    .B(_02356_),
    .Y(_02373_));
 sky130_fd_sc_hd__a21oi_1 _07192_ (.A1(_02372_),
    .A2(_02373_),
    .B1(net604),
    .Y(_00663_));
 sky130_fd_sc_hd__nand2_1 _07193_ (.A(net579),
    .B(net486),
    .Y(_02374_));
 sky130_fd_sc_hd__nand2_1 _07194_ (.A(\core.CPU_Dmem_value_a5[8][17] ),
    .B(net443),
    .Y(_02375_));
 sky130_fd_sc_hd__a21oi_1 _07195_ (.A1(_02374_),
    .A2(_02375_),
    .B1(net604),
    .Y(_00664_));
 sky130_fd_sc_hd__nand2_1 _07197_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net486),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_1 _07199_ (.A(\core.CPU_Dmem_value_a5[8][18] ),
    .B(_02356_),
    .Y(_02379_));
 sky130_fd_sc_hd__a21oi_1 _07200_ (.A1(_02377_),
    .A2(_02379_),
    .B1(net604),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _07201_ (.A(net578),
    .B(net487),
    .Y(_02380_));
 sky130_fd_sc_hd__nand2_1 _07202_ (.A(\core.CPU_Dmem_value_a5[8][19] ),
    .B(net443),
    .Y(_02381_));
 sky130_fd_sc_hd__a21oi_1 _07203_ (.A1(_02380_),
    .A2(_02381_),
    .B1(net600),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _07204_ (.A(net577),
    .B(net486),
    .Y(_02382_));
 sky130_fd_sc_hd__nand2_1 _07205_ (.A(\core.CPU_Dmem_value_a5[8][1] ),
    .B(net443),
    .Y(_02383_));
 sky130_fd_sc_hd__a21oi_1 _07207_ (.A1(_02382_),
    .A2(_02383_),
    .B1(net605),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _07208_ (.A(net576),
    .B(net487),
    .Y(_02385_));
 sky130_fd_sc_hd__nand2_1 _07209_ (.A(\core.CPU_Dmem_value_a5[8][20] ),
    .B(_02356_),
    .Y(_02386_));
 sky130_fd_sc_hd__a21oi_1 _07210_ (.A1(_02385_),
    .A2(_02386_),
    .B1(net601),
    .Y(_00668_));
 sky130_fd_sc_hd__nand2_1 _07211_ (.A(net575),
    .B(net487),
    .Y(_02387_));
 sky130_fd_sc_hd__nand2_1 _07212_ (.A(\core.CPU_Dmem_value_a5[8][21] ),
    .B(net443),
    .Y(_02388_));
 sky130_fd_sc_hd__a21oi_1 _07213_ (.A1(_02387_),
    .A2(_02388_),
    .B1(net601),
    .Y(_00669_));
 sky130_fd_sc_hd__nand2_1 _07214_ (.A(net574),
    .B(net487),
    .Y(_02389_));
 sky130_fd_sc_hd__nand2_1 _07215_ (.A(\core.CPU_Dmem_value_a5[8][22] ),
    .B(net443),
    .Y(_02390_));
 sky130_fd_sc_hd__a21oi_1 _07216_ (.A1(_02389_),
    .A2(_02390_),
    .B1(net601),
    .Y(_00670_));
 sky130_fd_sc_hd__nand2_1 _07217_ (.A(net573),
    .B(net487),
    .Y(_02391_));
 sky130_fd_sc_hd__nand2_1 _07218_ (.A(\core.CPU_Dmem_value_a5[8][23] ),
    .B(net443),
    .Y(_02392_));
 sky130_fd_sc_hd__a21oi_1 _07219_ (.A1(_02391_),
    .A2(_02392_),
    .B1(net601),
    .Y(_00671_));
 sky130_fd_sc_hd__nand2_1 _07220_ (.A(net572),
    .B(net487),
    .Y(_02393_));
 sky130_fd_sc_hd__nand2_1 _07221_ (.A(\core.CPU_Dmem_value_a5[8][24] ),
    .B(net443),
    .Y(_02394_));
 sky130_fd_sc_hd__a21oi_1 _07222_ (.A1(_02393_),
    .A2(_02394_),
    .B1(net601),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_1 _07223_ (.A(net571),
    .B(net487),
    .Y(_02395_));
 sky130_fd_sc_hd__nand2_1 _07224_ (.A(\core.CPU_Dmem_value_a5[8][25] ),
    .B(_02356_),
    .Y(_02396_));
 sky130_fd_sc_hd__a21oi_1 _07225_ (.A1(_02395_),
    .A2(_02396_),
    .B1(net601),
    .Y(_00673_));
 sky130_fd_sc_hd__nand2_1 _07226_ (.A(net570),
    .B(net486),
    .Y(_02397_));
 sky130_fd_sc_hd__nand2_1 _07227_ (.A(\core.CPU_Dmem_value_a5[8][26] ),
    .B(net443),
    .Y(_02398_));
 sky130_fd_sc_hd__a21oi_1 _07228_ (.A1(_02397_),
    .A2(_02398_),
    .B1(net603),
    .Y(_00674_));
 sky130_fd_sc_hd__nand2_1 _07230_ (.A(net569),
    .B(net486),
    .Y(_02400_));
 sky130_fd_sc_hd__nand2_1 _07232_ (.A(\core.CPU_Dmem_value_a5[8][27] ),
    .B(net443),
    .Y(_02402_));
 sky130_fd_sc_hd__a21oi_1 _07233_ (.A1(_02400_),
    .A2(_02402_),
    .B1(net604),
    .Y(_00675_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net486),
    .Y(_02403_));
 sky130_fd_sc_hd__nand2_1 _07235_ (.A(\core.CPU_Dmem_value_a5[8][28] ),
    .B(_02356_),
    .Y(_02404_));
 sky130_fd_sc_hd__a21oi_1 _07236_ (.A1(_02403_),
    .A2(_02404_),
    .B1(net603),
    .Y(_00676_));
 sky130_fd_sc_hd__nand2_1 _07237_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net487),
    .Y(_02405_));
 sky130_fd_sc_hd__nand2_1 _07238_ (.A(\core.CPU_Dmem_value_a5[8][29] ),
    .B(net443),
    .Y(_02406_));
 sky130_fd_sc_hd__a21oi_1 _07240_ (.A1(_02405_),
    .A2(_02406_),
    .B1(net599),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _07241_ (.A(net568),
    .B(net487),
    .Y(_02408_));
 sky130_fd_sc_hd__nand2_1 _07242_ (.A(\core.CPU_Dmem_value_a5[8][2] ),
    .B(net443),
    .Y(_02409_));
 sky130_fd_sc_hd__a21oi_1 _07243_ (.A1(_02408_),
    .A2(_02409_),
    .B1(net603),
    .Y(_00678_));
 sky130_fd_sc_hd__nand2_1 _07244_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net487),
    .Y(_02410_));
 sky130_fd_sc_hd__nand2_1 _07245_ (.A(\core.CPU_Dmem_value_a5[8][30] ),
    .B(_02356_),
    .Y(_02411_));
 sky130_fd_sc_hd__a21oi_1 _07246_ (.A1(_02410_),
    .A2(_02411_),
    .B1(net599),
    .Y(_00679_));
 sky130_fd_sc_hd__nand2_1 _07247_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net487),
    .Y(_02412_));
 sky130_fd_sc_hd__nand2_1 _07248_ (.A(\core.CPU_Dmem_value_a5[8][31] ),
    .B(net443),
    .Y(_02413_));
 sky130_fd_sc_hd__a21oi_1 _07249_ (.A1(_02412_),
    .A2(_02413_),
    .B1(net601),
    .Y(_00680_));
 sky130_fd_sc_hd__nand2_1 _07250_ (.A(\core.CPU_Dmem_value_a5[8][3] ),
    .B(_02356_),
    .Y(_02414_));
 sky130_fd_sc_hd__nand2_1 _07251_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net487),
    .Y(_02415_));
 sky130_fd_sc_hd__nand3b_1 _07252_ (.A_N(net599),
    .B(_02414_),
    .C(_02415_),
    .Y(_00681_));
 sky130_fd_sc_hd__nand2_1 _07253_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net486),
    .Y(_02416_));
 sky130_fd_sc_hd__nand2_1 _07254_ (.A(\core.CPU_Dmem_value_a5[8][4] ),
    .B(_02356_),
    .Y(_02417_));
 sky130_fd_sc_hd__a21oi_1 _07255_ (.A1(_02416_),
    .A2(_02417_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00682_));
 sky130_fd_sc_hd__nand2_1 _07256_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net486),
    .Y(_02418_));
 sky130_fd_sc_hd__nand2_1 _07257_ (.A(\core.CPU_Dmem_value_a5[8][5] ),
    .B(_02356_),
    .Y(_02419_));
 sky130_fd_sc_hd__a21oi_1 _07258_ (.A1(_02418_),
    .A2(_02419_),
    .B1(net605),
    .Y(_00683_));
 sky130_fd_sc_hd__nand2_1 _07259_ (.A(net567),
    .B(net487),
    .Y(_02420_));
 sky130_fd_sc_hd__nand2_1 _07260_ (.A(\core.CPU_Dmem_value_a5[8][6] ),
    .B(net443),
    .Y(_02421_));
 sky130_fd_sc_hd__a21oi_1 _07261_ (.A1(_02420_),
    .A2(_02421_),
    .B1(net599),
    .Y(_00684_));
 sky130_fd_sc_hd__nand2_1 _07262_ (.A(net566),
    .B(net487),
    .Y(_02422_));
 sky130_fd_sc_hd__nand2_1 _07263_ (.A(\core.CPU_Dmem_value_a5[8][7] ),
    .B(net443),
    .Y(_02423_));
 sky130_fd_sc_hd__a21oi_1 _07264_ (.A1(_02422_),
    .A2(_02423_),
    .B1(net599),
    .Y(_00685_));
 sky130_fd_sc_hd__nand2_1 _07265_ (.A(net565),
    .B(net487),
    .Y(_02424_));
 sky130_fd_sc_hd__nand2_1 _07266_ (.A(\core.CPU_Dmem_value_a5[8][8] ),
    .B(net443),
    .Y(_02425_));
 sky130_fd_sc_hd__a21oi_1 _07267_ (.A1(_02424_),
    .A2(_02425_),
    .B1(net601),
    .Y(_00686_));
 sky130_fd_sc_hd__nand2_1 _07268_ (.A(net564),
    .B(net487),
    .Y(_02426_));
 sky130_fd_sc_hd__nand2_1 _07269_ (.A(\core.CPU_Dmem_value_a5[8][9] ),
    .B(net443),
    .Y(_02427_));
 sky130_fd_sc_hd__a21oi_1 _07270_ (.A1(_02426_),
    .A2(_02427_),
    .B1(net603),
    .Y(_00687_));
 sky130_fd_sc_hd__nor2_4 _07271_ (.A(_01346_),
    .B(_01580_),
    .Y(_02428_));
 sky130_fd_sc_hd__nand2_2 _07273_ (.A(net560),
    .B(_02428_),
    .Y(_02430_));
 sky130_fd_sc_hd__nand2_1 _07275_ (.A(\core.CPU_Dmem_value_a5[9][0] ),
    .B(_02430_),
    .Y(_02432_));
 sky130_fd_sc_hd__nor3_2 _07276_ (.A(net561),
    .B(_01346_),
    .C(_01580_),
    .Y(_02433_));
 sky130_fd_sc_hd__nand2_1 _07278_ (.A(\core.CPU_dmem_wr_data_a4[0] ),
    .B(net482),
    .Y(_02435_));
 sky130_fd_sc_hd__nand3b_1 _07279_ (.A_N(\core.CPU_reset_a4 ),
    .B(_02432_),
    .C(_02435_),
    .Y(_00688_));
 sky130_fd_sc_hd__nand2_1 _07280_ (.A(net584),
    .B(net482),
    .Y(_02436_));
 sky130_fd_sc_hd__nand2_1 _07281_ (.A(\core.CPU_Dmem_value_a5[9][10] ),
    .B(net442),
    .Y(_02437_));
 sky130_fd_sc_hd__a21oi_1 _07283_ (.A1(_02436_),
    .A2(_02437_),
    .B1(net601),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _07284_ (.A(net583),
    .B(net482),
    .Y(_02439_));
 sky130_fd_sc_hd__nand2_1 _07285_ (.A(\core.CPU_Dmem_value_a5[9][11] ),
    .B(net442),
    .Y(_02440_));
 sky130_fd_sc_hd__a21oi_1 _07286_ (.A1(_02439_),
    .A2(_02440_),
    .B1(net601),
    .Y(_00690_));
 sky130_fd_sc_hd__nand2_1 _07287_ (.A(net582),
    .B(net482),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_1 _07288_ (.A(\core.CPU_Dmem_value_a5[9][12] ),
    .B(net442),
    .Y(_02442_));
 sky130_fd_sc_hd__a21oi_1 _07289_ (.A1(_02441_),
    .A2(_02442_),
    .B1(net600),
    .Y(_00691_));
 sky130_fd_sc_hd__nand2_1 _07290_ (.A(\core.CPU_dmem_wr_data_a4[13] ),
    .B(net482),
    .Y(_02443_));
 sky130_fd_sc_hd__nand2_1 _07291_ (.A(\core.CPU_Dmem_value_a5[9][13] ),
    .B(_02430_),
    .Y(_02444_));
 sky130_fd_sc_hd__a21oi_1 _07292_ (.A1(_02443_),
    .A2(_02444_),
    .B1(net604),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_1 _07293_ (.A(net581),
    .B(net482),
    .Y(_02445_));
 sky130_fd_sc_hd__nand2_1 _07294_ (.A(\core.CPU_Dmem_value_a5[9][14] ),
    .B(net442),
    .Y(_02446_));
 sky130_fd_sc_hd__a21oi_1 _07295_ (.A1(_02445_),
    .A2(_02446_),
    .B1(net602),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2_1 _07296_ (.A(net580),
    .B(net482),
    .Y(_02447_));
 sky130_fd_sc_hd__nand2_1 _07297_ (.A(\core.CPU_Dmem_value_a5[9][15] ),
    .B(net442),
    .Y(_02448_));
 sky130_fd_sc_hd__a21oi_1 _07298_ (.A1(_02447_),
    .A2(_02448_),
    .B1(net601),
    .Y(_00694_));
 sky130_fd_sc_hd__nand2_1 _07299_ (.A(\core.CPU_dmem_wr_data_a4[16] ),
    .B(net482),
    .Y(_02449_));
 sky130_fd_sc_hd__nand2_1 _07300_ (.A(\core.CPU_Dmem_value_a5[9][16] ),
    .B(_02430_),
    .Y(_02450_));
 sky130_fd_sc_hd__a21oi_1 _07301_ (.A1(_02449_),
    .A2(_02450_),
    .B1(net604),
    .Y(_00695_));
 sky130_fd_sc_hd__nand2_1 _07302_ (.A(net579),
    .B(net482),
    .Y(_02451_));
 sky130_fd_sc_hd__nand2_1 _07303_ (.A(\core.CPU_Dmem_value_a5[9][17] ),
    .B(_02430_),
    .Y(_02452_));
 sky130_fd_sc_hd__a21oi_1 _07304_ (.A1(_02451_),
    .A2(_02452_),
    .B1(net604),
    .Y(_00696_));
 sky130_fd_sc_hd__nand2_1 _07306_ (.A(\core.CPU_dmem_wr_data_a4[18] ),
    .B(net482),
    .Y(_02454_));
 sky130_fd_sc_hd__nand2_1 _07308_ (.A(\core.CPU_Dmem_value_a5[9][18] ),
    .B(_02430_),
    .Y(_02456_));
 sky130_fd_sc_hd__a21oi_1 _07309_ (.A1(_02454_),
    .A2(_02456_),
    .B1(net604),
    .Y(_00697_));
 sky130_fd_sc_hd__nand2_1 _07310_ (.A(net578),
    .B(net482),
    .Y(_02457_));
 sky130_fd_sc_hd__nand2_1 _07311_ (.A(\core.CPU_Dmem_value_a5[9][19] ),
    .B(net442),
    .Y(_02458_));
 sky130_fd_sc_hd__a21oi_1 _07312_ (.A1(_02457_),
    .A2(_02458_),
    .B1(net600),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _07313_ (.A(net577),
    .B(net482),
    .Y(_02459_));
 sky130_fd_sc_hd__nand2_1 _07314_ (.A(\core.CPU_Dmem_value_a5[9][1] ),
    .B(_02430_),
    .Y(_02460_));
 sky130_fd_sc_hd__a21oi_1 _07316_ (.A1(_02459_),
    .A2(_02460_),
    .B1(net605),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _07317_ (.A(net576),
    .B(net482),
    .Y(_02462_));
 sky130_fd_sc_hd__nand2_1 _07318_ (.A(\core.CPU_Dmem_value_a5[9][20] ),
    .B(net442),
    .Y(_02463_));
 sky130_fd_sc_hd__a21oi_1 _07319_ (.A1(_02462_),
    .A2(_02463_),
    .B1(net601),
    .Y(_00700_));
 sky130_fd_sc_hd__nand2_1 _07320_ (.A(net575),
    .B(net482),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2_1 _07321_ (.A(\core.CPU_Dmem_value_a5[9][21] ),
    .B(net442),
    .Y(_02465_));
 sky130_fd_sc_hd__a21oi_1 _07322_ (.A1(_02464_),
    .A2(_02465_),
    .B1(net601),
    .Y(_00701_));
 sky130_fd_sc_hd__nand2_1 _07323_ (.A(net574),
    .B(net482),
    .Y(_02466_));
 sky130_fd_sc_hd__nand2_1 _07324_ (.A(\core.CPU_Dmem_value_a5[9][22] ),
    .B(net442),
    .Y(_02467_));
 sky130_fd_sc_hd__a21oi_1 _07325_ (.A1(_02466_),
    .A2(_02467_),
    .B1(net601),
    .Y(_00702_));
 sky130_fd_sc_hd__nand2_1 _07326_ (.A(net573),
    .B(net482),
    .Y(_02468_));
 sky130_fd_sc_hd__nand2_1 _07327_ (.A(\core.CPU_Dmem_value_a5[9][23] ),
    .B(net442),
    .Y(_02469_));
 sky130_fd_sc_hd__a21oi_1 _07328_ (.A1(_02468_),
    .A2(_02469_),
    .B1(net601),
    .Y(_00703_));
 sky130_fd_sc_hd__nand2_1 _07329_ (.A(net572),
    .B(net482),
    .Y(_02470_));
 sky130_fd_sc_hd__nand2_1 _07330_ (.A(\core.CPU_Dmem_value_a5[9][24] ),
    .B(net442),
    .Y(_02471_));
 sky130_fd_sc_hd__a21oi_1 _07331_ (.A1(_02470_),
    .A2(_02471_),
    .B1(net601),
    .Y(_00704_));
 sky130_fd_sc_hd__nand2_1 _07332_ (.A(net571),
    .B(net482),
    .Y(_02472_));
 sky130_fd_sc_hd__nand2_1 _07333_ (.A(\core.CPU_Dmem_value_a5[9][25] ),
    .B(net442),
    .Y(_02473_));
 sky130_fd_sc_hd__a21oi_1 _07334_ (.A1(_02472_),
    .A2(_02473_),
    .B1(net601),
    .Y(_00705_));
 sky130_fd_sc_hd__nand2_1 _07335_ (.A(net570),
    .B(net482),
    .Y(_02474_));
 sky130_fd_sc_hd__nand2_1 _07336_ (.A(\core.CPU_Dmem_value_a5[9][26] ),
    .B(_02430_),
    .Y(_02475_));
 sky130_fd_sc_hd__a21oi_1 _07337_ (.A1(_02474_),
    .A2(_02475_),
    .B1(net603),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_1 _07339_ (.A(net569),
    .B(net482),
    .Y(_02477_));
 sky130_fd_sc_hd__nand2_1 _07341_ (.A(\core.CPU_Dmem_value_a5[9][27] ),
    .B(_02430_),
    .Y(_02479_));
 sky130_fd_sc_hd__a21oi_1 _07342_ (.A1(_02477_),
    .A2(_02479_),
    .B1(net604),
    .Y(_00707_));
 sky130_fd_sc_hd__nand2_1 _07343_ (.A(\core.CPU_dmem_wr_data_a4[28] ),
    .B(net482),
    .Y(_02480_));
 sky130_fd_sc_hd__nand2_1 _07344_ (.A(\core.CPU_Dmem_value_a5[9][28] ),
    .B(_02430_),
    .Y(_02481_));
 sky130_fd_sc_hd__a21oi_1 _07345_ (.A1(_02480_),
    .A2(_02481_),
    .B1(net603),
    .Y(_00708_));
 sky130_fd_sc_hd__nand2_1 _07346_ (.A(\core.CPU_dmem_wr_data_a4[29] ),
    .B(net482),
    .Y(_02482_));
 sky130_fd_sc_hd__nand2_1 _07347_ (.A(\core.CPU_Dmem_value_a5[9][29] ),
    .B(net442),
    .Y(_02483_));
 sky130_fd_sc_hd__a21oi_1 _07349_ (.A1(_02482_),
    .A2(_02483_),
    .B1(net602),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _07350_ (.A(net568),
    .B(net482),
    .Y(_02485_));
 sky130_fd_sc_hd__nand2_1 _07351_ (.A(\core.CPU_Dmem_value_a5[9][2] ),
    .B(net442),
    .Y(_02486_));
 sky130_fd_sc_hd__a21oi_1 _07352_ (.A1(_02485_),
    .A2(_02486_),
    .B1(net603),
    .Y(_00710_));
 sky130_fd_sc_hd__nand2_1 _07353_ (.A(\core.CPU_dmem_wr_data_a4[30] ),
    .B(net482),
    .Y(_02487_));
 sky130_fd_sc_hd__nand2_1 _07354_ (.A(\core.CPU_Dmem_value_a5[9][30] ),
    .B(net442),
    .Y(_02488_));
 sky130_fd_sc_hd__a21oi_1 _07355_ (.A1(_02487_),
    .A2(_02488_),
    .B1(net602),
    .Y(_00711_));
 sky130_fd_sc_hd__nand2_1 _07356_ (.A(\core.CPU_dmem_wr_data_a4[31] ),
    .B(net482),
    .Y(_02489_));
 sky130_fd_sc_hd__nand2_1 _07357_ (.A(\core.CPU_Dmem_value_a5[9][31] ),
    .B(net442),
    .Y(_02490_));
 sky130_fd_sc_hd__a21oi_1 _07358_ (.A1(_02489_),
    .A2(_02490_),
    .B1(net601),
    .Y(_00712_));
 sky130_fd_sc_hd__nand2_1 _07359_ (.A(\core.CPU_Dmem_value_a5[9][3] ),
    .B(net442),
    .Y(_02491_));
 sky130_fd_sc_hd__nand2_1 _07360_ (.A(\core.CPU_dmem_wr_data_a4[3] ),
    .B(net482),
    .Y(_02492_));
 sky130_fd_sc_hd__nand3b_1 _07361_ (.A_N(net602),
    .B(_02491_),
    .C(_02492_),
    .Y(_00713_));
 sky130_fd_sc_hd__nand2_1 _07362_ (.A(\core.CPU_dmem_wr_data_a4[4] ),
    .B(net482),
    .Y(_02493_));
 sky130_fd_sc_hd__nand2_1 _07363_ (.A(\core.CPU_Dmem_value_a5[9][4] ),
    .B(net442),
    .Y(_02494_));
 sky130_fd_sc_hd__a21oi_1 _07364_ (.A1(_02493_),
    .A2(_02494_),
    .B1(\core.CPU_reset_a4 ),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2_1 _07365_ (.A(\core.CPU_dmem_wr_data_a4[5] ),
    .B(net482),
    .Y(_02495_));
 sky130_fd_sc_hd__nand2_1 _07366_ (.A(\core.CPU_Dmem_value_a5[9][5] ),
    .B(_02430_),
    .Y(_02496_));
 sky130_fd_sc_hd__a21oi_1 _07367_ (.A1(_02495_),
    .A2(_02496_),
    .B1(net604),
    .Y(_00715_));
 sky130_fd_sc_hd__nand2_1 _07368_ (.A(net567),
    .B(net482),
    .Y(_02497_));
 sky130_fd_sc_hd__nand2_1 _07369_ (.A(\core.CPU_Dmem_value_a5[9][6] ),
    .B(net442),
    .Y(_02498_));
 sky130_fd_sc_hd__a21oi_1 _07370_ (.A1(_02497_),
    .A2(_02498_),
    .B1(net602),
    .Y(_00716_));
 sky130_fd_sc_hd__nand2_1 _07371_ (.A(net566),
    .B(net482),
    .Y(_02499_));
 sky130_fd_sc_hd__nand2_1 _07372_ (.A(\core.CPU_Dmem_value_a5[9][7] ),
    .B(net442),
    .Y(_02500_));
 sky130_fd_sc_hd__a21oi_1 _07373_ (.A1(_02499_),
    .A2(_02500_),
    .B1(net602),
    .Y(_00717_));
 sky130_fd_sc_hd__nand2_1 _07374_ (.A(net565),
    .B(net482),
    .Y(_02501_));
 sky130_fd_sc_hd__nand2_1 _07375_ (.A(\core.CPU_Dmem_value_a5[9][8] ),
    .B(net442),
    .Y(_02502_));
 sky130_fd_sc_hd__a21oi_1 _07376_ (.A1(_02501_),
    .A2(_02502_),
    .B1(net601),
    .Y(_00718_));
 sky130_fd_sc_hd__nand2_1 _07377_ (.A(net564),
    .B(net482),
    .Y(_02503_));
 sky130_fd_sc_hd__nand2_1 _07378_ (.A(\core.CPU_Dmem_value_a5[9][9] ),
    .B(net442),
    .Y(_02504_));
 sky130_fd_sc_hd__a21oi_1 _07379_ (.A1(_02503_),
    .A2(_02504_),
    .B1(net603),
    .Y(_00719_));
 sky130_fd_sc_hd__nor2b_1 _07383_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][0] ),
    .Y(_00720_));
 sky130_fd_sc_hd__nor2b_1 _07385_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][10] ),
    .Y(_00721_));
 sky130_fd_sc_hd__nor2b_1 _07386_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][11] ),
    .Y(_00722_));
 sky130_fd_sc_hd__nor2b_1 _07387_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][12] ),
    .Y(_00723_));
 sky130_fd_sc_hd__nor2b_1 _07388_ (.A(\core.CPU_reset_a3 ),
    .B_N(\core.CPU_Xreg_value_a4[0][13] ),
    .Y(_00724_));
 sky130_fd_sc_hd__nor2b_1 _07389_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][14] ),
    .Y(_00725_));
 sky130_fd_sc_hd__nor2b_1 _07390_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][15] ),
    .Y(_00726_));
 sky130_fd_sc_hd__nor2b_1 _07391_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][16] ),
    .Y(_00727_));
 sky130_fd_sc_hd__nor2b_1 _07392_ (.A(\core.CPU_reset_a3 ),
    .B_N(\core.CPU_Xreg_value_a4[0][17] ),
    .Y(_00728_));
 sky130_fd_sc_hd__nor2b_1 _07393_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][18] ),
    .Y(_00729_));
 sky130_fd_sc_hd__nor2b_1 _07394_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][19] ),
    .Y(_00730_));
 sky130_fd_sc_hd__nor2b_1 _07396_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][1] ),
    .Y(_00731_));
 sky130_fd_sc_hd__nor2b_1 _07397_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][20] ),
    .Y(_00732_));
 sky130_fd_sc_hd__nor2b_1 _07398_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][21] ),
    .Y(_00733_));
 sky130_fd_sc_hd__nor2b_1 _07399_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][22] ),
    .Y(_00734_));
 sky130_fd_sc_hd__nor2b_1 _07400_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][23] ),
    .Y(_00735_));
 sky130_fd_sc_hd__nor2b_1 _07401_ (.A(\core.CPU_reset_a3 ),
    .B_N(\core.CPU_Xreg_value_a4[0][24] ),
    .Y(_00736_));
 sky130_fd_sc_hd__nor2b_1 _07402_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][25] ),
    .Y(_00737_));
 sky130_fd_sc_hd__nor2b_1 _07403_ (.A(\core.CPU_reset_a3 ),
    .B_N(\core.CPU_Xreg_value_a4[0][26] ),
    .Y(_00738_));
 sky130_fd_sc_hd__nor2b_1 _07404_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][27] ),
    .Y(_00739_));
 sky130_fd_sc_hd__nor2b_1 _07405_ (.A(\core.CPU_reset_a3 ),
    .B_N(\core.CPU_Xreg_value_a4[0][28] ),
    .Y(_00740_));
 sky130_fd_sc_hd__nor2b_1 _07407_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][29] ),
    .Y(_00741_));
 sky130_fd_sc_hd__nor2b_1 _07408_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][2] ),
    .Y(_00742_));
 sky130_fd_sc_hd__nor2b_1 _07409_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][30] ),
    .Y(_00743_));
 sky130_fd_sc_hd__nor2b_1 _07410_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][31] ),
    .Y(_00744_));
 sky130_fd_sc_hd__nor2b_1 _07411_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][3] ),
    .Y(_00745_));
 sky130_fd_sc_hd__nor2b_1 _07412_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][4] ),
    .Y(_00746_));
 sky130_fd_sc_hd__nor2b_1 _07413_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][5] ),
    .Y(_00747_));
 sky130_fd_sc_hd__nor2b_1 _07414_ (.A(net607),
    .B_N(\core.CPU_Xreg_value_a4[0][6] ),
    .Y(_00748_));
 sky130_fd_sc_hd__nor2b_1 _07415_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][7] ),
    .Y(_00749_));
 sky130_fd_sc_hd__nor2b_1 _07416_ (.A(net606),
    .B_N(\core.CPU_Xreg_value_a4[0][8] ),
    .Y(_00750_));
 sky130_fd_sc_hd__nor2b_1 _07418_ (.A(\core.CPU_reset_a3 ),
    .B_N(\core.CPU_Xreg_value_a4[0][9] ),
    .Y(_00751_));
 sky130_fd_sc_hd__inv_1 _07419_ (.A(\core.CPU_is_addi_a3 ),
    .Y(_02512_));
 sky130_fd_sc_hd__nor2_1 _07424_ (.A(net609),
    .B(net612),
    .Y(_02517_));
 sky130_fd_sc_hd__nor2_1 _07428_ (.A(net610),
    .B(_00038_),
    .Y(_02521_));
 sky130_fd_sc_hd__or3b_2 _07430_ (.A(\core.CPU_imm_a3[4] ),
    .B(\core.CPU_imm_a3[5] ),
    .C_N(net610),
    .X(_02523_));
 sky130_fd_sc_hd__or3b_1 _07431_ (.A(net610),
    .B(\core.CPU_src2_value_a3[4] ),
    .C_N(\core.CPU_is_sll_a3 ),
    .X(_02524_));
 sky130_fd_sc_hd__and2_1 _07432_ (.A(_02523_),
    .B(_02524_),
    .X(_02525_));
 sky130_fd_sc_hd__nand2_1 _07434_ (.A(net610),
    .B(\core.CPU_imm_a3[3] ),
    .Y(_02527_));
 sky130_fd_sc_hd__o21ai_2 _07435_ (.A1(net610),
    .A2(_00044_),
    .B1(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__nor3_1 _07437_ (.A(net481),
    .B(_02525_),
    .C(net480),
    .Y(_02530_));
 sky130_fd_sc_hd__or3b_2 _07438_ (.A(\core.CPU_imm_a3[0] ),
    .B(\core.CPU_imm_a3[1] ),
    .C_N(net610),
    .X(_02531_));
 sky130_fd_sc_hd__or3_1 _07439_ (.A(\core.CPU_src2_value_a3[0] ),
    .B(net610),
    .C(\core.CPU_src2_value_a3[1] ),
    .X(_02532_));
 sky130_fd_sc_hd__a21oi_1 _07440_ (.A1(_02531_),
    .A2(_02532_),
    .B1(_00021_),
    .Y(_02533_));
 sky130_fd_sc_hd__nand3_1 _07441_ (.A(_02517_),
    .B(net441),
    .C(net479),
    .Y(_02534_));
 sky130_fd_sc_hd__o21ai_0 _07442_ (.A1(_00022_),
    .A2(_02517_),
    .B1(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__inv_1 _07443_ (.A(\core.CPU_is_sub_a3 ),
    .Y(_02536_));
 sky130_fd_sc_hd__inv_1 _07444_ (.A(net612),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2_1 _07446_ (.A(net556),
    .B(net555),
    .Y(_02539_));
 sky130_fd_sc_hd__or2_2 _07447_ (.A(net610),
    .B(\core.CPU_is_sll_a3 ),
    .X(_02540_));
 sky130_fd_sc_hd__o21ai_0 _07449_ (.A1(_02539_),
    .A2(_02540_),
    .B1(net557),
    .Y(_02542_));
 sky130_fd_sc_hd__a22oi_1 _07450_ (.A1(net557),
    .A2(_02535_),
    .B1(_02542_),
    .B2(_00031_),
    .Y(_02543_));
 sky130_fd_sc_hd__nor2_1 _07451_ (.A(\core.CPU_dmem_rd_data_a5[0] ),
    .B(net536),
    .Y(_02544_));
 sky130_fd_sc_hd__a21oi_1 _07452_ (.A1(net535),
    .A2(net394),
    .B1(net440),
    .Y(_02545_));
 sky130_fd_sc_hd__nand2b_1 _07453_ (.A_N(\core.CPU_rd_a5[4] ),
    .B(\core.CPU_rd_a5[3] ),
    .Y(_02546_));
 sky130_fd_sc_hd__inv_1 _07455_ (.A(\core.CPU_rd_a3[4] ),
    .Y(_02548_));
 sky130_fd_sc_hd__nand3_1 _07456_ (.A(\core.CPU_rd_a3[3] ),
    .B(_02548_),
    .C(net535),
    .Y(_02549_));
 sky130_fd_sc_hd__o21a_1 _07457_ (.A1(net535),
    .A2(_02546_),
    .B1(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__nor3b_1 _07458_ (.A(_01114_),
    .B(\core.CPU_rd_a3[0] ),
    .C_N(\core.CPU_rd_a3[1] ),
    .Y(_02551_));
 sky130_fd_sc_hd__nor3b_1 _07459_ (.A(\core.CPU_rd_a5[0] ),
    .B(net535),
    .C_N(\core.CPU_rd_a5[1] ),
    .Y(_02552_));
 sky130_fd_sc_hd__nor2_1 _07460_ (.A(\core.CPU_rd_a3[0] ),
    .B(\core.CPU_rd_a3[1] ),
    .Y(_02553_));
 sky130_fd_sc_hd__nor2_1 _07461_ (.A(\core.CPU_rd_a3[3] ),
    .B(\core.CPU_rd_a3[4] ),
    .Y(_02554_));
 sky130_fd_sc_hd__nand2_1 _07462_ (.A(_02553_),
    .B(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__a31o_2 _07463_ (.A1(\core.CPU_rd_valid_a3 ),
    .A2(net535),
    .A3(_02555_),
    .B1(\core.CPU_valid_load_a5 ),
    .X(_02556_));
 sky130_fd_sc_hd__o21ai_1 _07464_ (.A1(_02551_),
    .A2(_02552_),
    .B1(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__nor2_2 _07465_ (.A(_02550_),
    .B(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__nand2_1 _07467_ (.A(_02545_),
    .B(_02558_),
    .Y(_02560_));
 sky130_fd_sc_hd__o21ai_0 _07468_ (.A1(net535),
    .A2(_02546_),
    .B1(_02549_),
    .Y(_02561_));
 sky130_fd_sc_hd__o21a_1 _07469_ (.A1(_02551_),
    .A2(_02552_),
    .B1(_02556_),
    .X(_02562_));
 sky130_fd_sc_hd__nand2_2 _07470_ (.A(_02561_),
    .B(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__nand2_1 _07473_ (.A(\core.CPU_Xreg_value_a4[10][0] ),
    .B(net428),
    .Y(_02566_));
 sky130_fd_sc_hd__a21oi_1 _07475_ (.A1(_02560_),
    .A2(_02566_),
    .B1(net607),
    .Y(_00752_));
 sky130_fd_sc_hd__mux2i_4 _07478_ (.A0(\core.CPU_src2_value_a3[0] ),
    .A1(\core.CPU_imm_a3[0] ),
    .S(net610),
    .Y(_02570_));
 sky130_fd_sc_hd__mux2i_1 _07480_ (.A0(\core.CPU_src1_value_a3[5] ),
    .A1(\core.CPU_src1_value_a3[6] ),
    .S(net554),
    .Y(_02572_));
 sky130_fd_sc_hd__mux2i_1 _07481_ (.A0(\core.CPU_src1_value_a3[3] ),
    .A1(\core.CPU_src1_value_a3[4] ),
    .S(net554),
    .Y(_02573_));
 sky130_fd_sc_hd__mux2i_1 _07483_ (.A0(\core.CPU_src1_value_a3[9] ),
    .A1(\core.CPU_src1_value_a3[10] ),
    .S(net554),
    .Y(_02575_));
 sky130_fd_sc_hd__mux2i_1 _07484_ (.A0(\core.CPU_src1_value_a3[7] ),
    .A1(\core.CPU_src1_value_a3[8] ),
    .S(net554),
    .Y(_02576_));
 sky130_fd_sc_hd__mux2_2 _07485_ (.A0(\core.CPU_src2_value_a3[1] ),
    .A1(\core.CPU_imm_a3[1] ),
    .S(net610),
    .X(_02577_));
 sky130_fd_sc_hd__nand2b_1 _07486_ (.A_N(net610),
    .B(\core.CPU_src2_value_a3[2] ),
    .Y(_02578_));
 sky130_fd_sc_hd__mux4_2 _07488_ (.A0(_02572_),
    .A1(_02573_),
    .A2(_02575_),
    .A3(_02576_),
    .S0(_02577_),
    .S1(net553),
    .X(_02580_));
 sky130_fd_sc_hd__inv_1 _07489_ (.A(\core.CPU_imm_a3[0] ),
    .Y(_02581_));
 sky130_fd_sc_hd__nor2_1 _07490_ (.A(\core.CPU_src2_value_a3[0] ),
    .B(net610),
    .Y(_02582_));
 sky130_fd_sc_hd__a32oi_1 _07491_ (.A1(_02581_),
    .A2(net610),
    .A3(\core.CPU_imm_a3[1] ),
    .B1(_02582_),
    .B2(\core.CPU_src2_value_a3[1] ),
    .Y(_02583_));
 sky130_fd_sc_hd__mux2i_1 _07493_ (.A0(\core.CPU_src1_value_a3[1] ),
    .A1(\core.CPU_src1_value_a3[2] ),
    .S(_02570_),
    .Y(_02585_));
 sky130_fd_sc_hd__o22ai_1 _07494_ (.A1(_00021_),
    .A2(_02583_),
    .B1(_02585_),
    .B2(_02577_),
    .Y(_02586_));
 sky130_fd_sc_hd__o21a_1 _07495_ (.A1(net610),
    .A2(_00044_),
    .B1(_02527_),
    .X(_02587_));
 sky130_fd_sc_hd__nor2_1 _07496_ (.A(net481),
    .B(net478),
    .Y(_02588_));
 sky130_fd_sc_hd__a2bb2oi_1 _07497_ (.A1_N(net480),
    .A2_N(_02580_),
    .B1(_02586_),
    .B2(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__o21ai_0 _07498_ (.A1(_02525_),
    .A2(_02589_),
    .B1(_02517_),
    .Y(_02590_));
 sky130_fd_sc_hd__inv_1 _07500_ (.A(_00080_),
    .Y(_02592_));
 sky130_fd_sc_hd__a21oi_1 _07501_ (.A1(_02592_),
    .A2(_00077_),
    .B1(_00081_),
    .Y(_02593_));
 sky130_fd_sc_hd__nor2b_1 _07502_ (.A(_00040_),
    .B_N(_00008_),
    .Y(_02594_));
 sky130_fd_sc_hd__or2_2 _07503_ (.A(_00041_),
    .B(_00047_),
    .X(_02595_));
 sky130_fd_sc_hd__nand2b_1 _07504_ (.A_N(_00047_),
    .B(_00046_),
    .Y(_02596_));
 sky130_fd_sc_hd__nor2_1 _07505_ (.A(_00052_),
    .B(_00056_),
    .Y(_02597_));
 sky130_fd_sc_hd__o211a_1 _07506_ (.A1(_02594_),
    .A2(_02595_),
    .B1(_02596_),
    .C1(_02597_),
    .X(_02598_));
 sky130_fd_sc_hd__inv_1 _07507_ (.A(_00053_),
    .Y(_02599_));
 sky130_fd_sc_hd__inv_1 _07508_ (.A(_00057_),
    .Y(_02600_));
 sky130_fd_sc_hd__inv_1 _07509_ (.A(_00071_),
    .Y(_02601_));
 sky130_fd_sc_hd__nand2b_1 _07510_ (.A_N(_00070_),
    .B(_00063_),
    .Y(_02602_));
 sky130_fd_sc_hd__o2111ai_1 _07511_ (.A1(_02599_),
    .A2(_00056_),
    .B1(_02600_),
    .C1(_02601_),
    .D1(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__nor3b_1 _07512_ (.A(_00063_),
    .B(_00071_),
    .C_N(_00062_),
    .Y(_02604_));
 sky130_fd_sc_hd__a2111oi_0 _07513_ (.A1(_00070_),
    .A2(_02601_),
    .B1(_00076_),
    .C1(_00080_),
    .D1(_02604_),
    .Y(_02605_));
 sky130_fd_sc_hd__o21ai_0 _07514_ (.A1(_02598_),
    .A2(_02603_),
    .B1(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__nand2_1 _07515_ (.A(_02593_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__xnor2_1 _07516_ (.A(_00086_),
    .B(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(net609),
    .B(net555),
    .Y(_02609_));
 sky130_fd_sc_hd__inv_1 _07518_ (.A(_00086_),
    .Y(_02610_));
 sky130_fd_sc_hd__nor2b_1 _07519_ (.A(_00005_),
    .B_N(_00040_),
    .Y(_02611_));
 sky130_fd_sc_hd__o21a_1 _07520_ (.A1(_00046_),
    .A2(_00045_),
    .B1(_00052_),
    .X(_02612_));
 sky130_fd_sc_hd__o31a_1 _07521_ (.A1(_00039_),
    .A2(_00045_),
    .A3(_02611_),
    .B1(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__nand2_1 _07522_ (.A(_00056_),
    .B(_00062_),
    .Y(_02614_));
 sky130_fd_sc_hd__nor2_1 _07523_ (.A(_01146_),
    .B(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__o21ai_0 _07524_ (.A1(_00051_),
    .A2(_02613_),
    .B1(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_1 _07525_ (.A(_00062_),
    .B(_00055_),
    .Y(_02617_));
 sky130_fd_sc_hd__nor2_1 _07526_ (.A(_01146_),
    .B(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__nand2_1 _07527_ (.A(_00076_),
    .B(_00080_),
    .Y(_02619_));
 sky130_fd_sc_hd__a21oi_1 _07528_ (.A1(_00070_),
    .A2(_00061_),
    .B1(_00069_),
    .Y(_02620_));
 sky130_fd_sc_hd__a21oi_1 _07529_ (.A1(_00080_),
    .A2(_00075_),
    .B1(_00079_),
    .Y(_02621_));
 sky130_fd_sc_hd__o21ai_0 _07530_ (.A1(_02619_),
    .A2(_02620_),
    .B1(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__nor2_1 _07531_ (.A(_02618_),
    .B(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__nand2_1 _07532_ (.A(_02616_),
    .B(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__xnor2_1 _07533_ (.A(_02610_),
    .B(_02624_),
    .Y(_02625_));
 sky130_fd_sc_hd__o22ai_1 _07534_ (.A1(net555),
    .A2(_02608_),
    .B1(_02609_),
    .B2(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__nor2_1 _07535_ (.A(net611),
    .B(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__a21oi_1 _07536_ (.A1(_00065_),
    .A2(_00066_),
    .B1(_00064_),
    .Y(_02628_));
 sky130_fd_sc_hd__inv_1 _07537_ (.A(_00058_),
    .Y(_02629_));
 sky130_fd_sc_hd__o21ai_0 _07538_ (.A1(_00049_),
    .A2(_00048_),
    .B1(_00059_),
    .Y(_02630_));
 sky130_fd_sc_hd__a31oi_1 _07539_ (.A1(_00001_),
    .A2(\core.CPU_src1_value_a3[2] ),
    .A3(_00043_),
    .B1(_00042_),
    .Y(_02631_));
 sky130_fd_sc_hd__nor2_1 _07540_ (.A(_00048_),
    .B(_00058_),
    .Y(_02632_));
 sky130_fd_sc_hd__nand2_1 _07541_ (.A(_00067_),
    .B(_00065_),
    .Y(_02633_));
 sky130_fd_sc_hd__a221o_1 _07542_ (.A1(_02629_),
    .A2(_02630_),
    .B1(_02631_),
    .B2(_02632_),
    .C1(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__nand2_1 _07543_ (.A(_02628_),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__a21o_1 _07544_ (.A1(_00073_),
    .A2(_02635_),
    .B1(_00072_),
    .X(_02636_));
 sky130_fd_sc_hd__a21oi_1 _07545_ (.A1(_00083_),
    .A2(_02636_),
    .B1(_00082_),
    .Y(_02637_));
 sky130_fd_sc_hd__xnor2_1 _07546_ (.A(_00089_),
    .B(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__o21ai_0 _07547_ (.A1(_02540_),
    .A2(_02626_),
    .B1(net557),
    .Y(_02639_));
 sky130_fd_sc_hd__a22oi_1 _07548_ (.A1(_02590_),
    .A2(_02627_),
    .B1(_02638_),
    .B2(_02639_),
    .Y(_02640_));
 sky130_fd_sc_hd__nor2_1 _07549_ (.A(\core.CPU_dmem_rd_data_a5[10] ),
    .B(net536),
    .Y(_02641_));
 sky130_fd_sc_hd__a211o_1 _07550_ (.A1(net536),
    .A2(_02640_),
    .B1(_02641_),
    .C1(\core.CPU_reset_a3 ),
    .X(_02642_));
 sky130_fd_sc_hd__inv_8 _07552_ (.A(\core.CPU_reset_a3 ),
    .Y(_02644_));
 sky130_fd_sc_hd__nand3_1 _07557_ (.A(\core.CPU_Xreg_value_a4[10][10] ),
    .B(net550),
    .C(net428),
    .Y(_02649_));
 sky130_fd_sc_hd__o21ai_0 _07558_ (.A1(net428),
    .A2(net348),
    .B1(_02649_),
    .Y(_00753_));
 sky130_fd_sc_hd__nor2_1 _07559_ (.A(\core.CPU_dmem_rd_data_a5[11] ),
    .B(net536),
    .Y(_02650_));
 sky130_fd_sc_hd__a21oi_1 _07560_ (.A1(_00089_),
    .A2(_00082_),
    .B1(_00088_),
    .Y(_02651_));
 sky130_fd_sc_hd__a21oi_1 _07561_ (.A1(_00073_),
    .A2(_00064_),
    .B1(_00072_),
    .Y(_02652_));
 sky130_fd_sc_hd__nand2_1 _07562_ (.A(_02651_),
    .B(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__a211oi_1 _07563_ (.A1(_00000_),
    .A2(_00033_),
    .B1(_00032_),
    .C1(_00042_),
    .Y(_02654_));
 sky130_fd_sc_hd__a21oi_1 _07564_ (.A1(\core.CPU_src1_value_a3[2] ),
    .A2(_00043_),
    .B1(_00042_),
    .Y(_02655_));
 sky130_fd_sc_hd__nand3_1 _07565_ (.A(_00059_),
    .B(_00067_),
    .C(_00049_),
    .Y(_02656_));
 sky130_fd_sc_hd__nor3_1 _07566_ (.A(_02654_),
    .B(_02655_),
    .C(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__nand3_1 _07567_ (.A(_00059_),
    .B(_00067_),
    .C(_00048_),
    .Y(_02658_));
 sky130_fd_sc_hd__a21oi_1 _07568_ (.A1(_00067_),
    .A2(_00058_),
    .B1(_00066_),
    .Y(_02659_));
 sky130_fd_sc_hd__nand2_1 _07569_ (.A(_02658_),
    .B(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__nand2_1 _07570_ (.A(_00065_),
    .B(_00073_),
    .Y(_02661_));
 sky130_fd_sc_hd__o21ai_0 _07571_ (.A1(_00083_),
    .A2(_00082_),
    .B1(_00089_),
    .Y(_02662_));
 sky130_fd_sc_hd__inv_1 _07572_ (.A(_00088_),
    .Y(_02663_));
 sky130_fd_sc_hd__a32oi_1 _07573_ (.A1(_02651_),
    .A2(_02652_),
    .A3(_02661_),
    .B1(_02662_),
    .B2(_02663_),
    .Y(_02664_));
 sky130_fd_sc_hd__o31ai_2 _07574_ (.A1(_02653_),
    .A2(_02657_),
    .A3(_02660_),
    .B1(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__xor2_1 _07575_ (.A(_00095_),
    .B(net435),
    .X(_02666_));
 sky130_fd_sc_hd__nand2_1 _07576_ (.A(_02523_),
    .B(_02524_),
    .Y(_02667_));
 sky130_fd_sc_hd__mux2i_1 _07577_ (.A0(\core.CPU_src1_value_a3[2] ),
    .A1(\core.CPU_src1_value_a3[0] ),
    .S(_02577_),
    .Y(_02668_));
 sky130_fd_sc_hd__mux2i_1 _07578_ (.A0(\core.CPU_src1_value_a3[3] ),
    .A1(\core.CPU_src1_value_a3[1] ),
    .S(_02577_),
    .Y(_02669_));
 sky130_fd_sc_hd__mux2i_1 _07579_ (.A0(_02668_),
    .A1(_02669_),
    .S(net554),
    .Y(_02670_));
 sky130_fd_sc_hd__mux2i_4 _07580_ (.A0(\core.CPU_src2_value_a3[1] ),
    .A1(\core.CPU_imm_a3[1] ),
    .S(net610),
    .Y(_02671_));
 sky130_fd_sc_hd__mux4_2 _07581_ (.A0(\core.CPU_src1_value_a3[8] ),
    .A1(\core.CPU_src1_value_a3[9] ),
    .A2(\core.CPU_src1_value_a3[10] ),
    .A3(\core.CPU_src1_value_a3[11] ),
    .S0(net554),
    .S1(net548),
    .X(_02672_));
 sky130_fd_sc_hd__and2_1 _07582_ (.A(net478),
    .B(_02672_),
    .X(_02673_));
 sky130_fd_sc_hd__a211o_1 _07583_ (.A1(net480),
    .A2(_02670_),
    .B1(_02673_),
    .C1(net481),
    .X(_02674_));
 sky130_fd_sc_hd__mux2i_1 _07584_ (.A0(\core.CPU_src1_value_a3[4] ),
    .A1(\core.CPU_src1_value_a3[6] ),
    .S(net548),
    .Y(_02675_));
 sky130_fd_sc_hd__mux2i_1 _07585_ (.A0(\core.CPU_src1_value_a3[5] ),
    .A1(\core.CPU_src1_value_a3[7] ),
    .S(net548),
    .Y(_02676_));
 sky130_fd_sc_hd__mux2_2 _07586_ (.A0(_02675_),
    .A1(_02676_),
    .S(net554),
    .X(_02677_));
 sky130_fd_sc_hd__o21ai_0 _07587_ (.A1(net480),
    .A2(_02677_),
    .B1(net481),
    .Y(_02678_));
 sky130_fd_sc_hd__a31oi_1 _07588_ (.A1(_02667_),
    .A2(_02674_),
    .A3(_02678_),
    .B1(_02539_),
    .Y(_02679_));
 sky130_fd_sc_hd__o22ai_1 _07589_ (.A1(_02540_),
    .A2(_02666_),
    .B1(_02679_),
    .B2(net611),
    .Y(_02680_));
 sky130_fd_sc_hd__nor2_1 _07590_ (.A(net556),
    .B(net612),
    .Y(_02681_));
 sky130_fd_sc_hd__inv_1 _07591_ (.A(_00092_),
    .Y(_02682_));
 sky130_fd_sc_hd__nand2_1 _07592_ (.A(_00080_),
    .B(_00086_),
    .Y(_02683_));
 sky130_fd_sc_hd__a21oi_1 _07593_ (.A1(_00076_),
    .A2(_00069_),
    .B1(_00075_),
    .Y(_02684_));
 sky130_fd_sc_hd__a21oi_1 _07594_ (.A1(_00086_),
    .A2(_00079_),
    .B1(_00085_),
    .Y(_02685_));
 sky130_fd_sc_hd__o21ai_0 _07595_ (.A1(_02683_),
    .A2(_02684_),
    .B1(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hd__nand2b_1 _07596_ (.A_N(_00004_),
    .B(_00034_),
    .Y(_02687_));
 sky130_fd_sc_hd__nor2_1 _07597_ (.A(_00036_),
    .B(_00039_),
    .Y(_02688_));
 sky130_fd_sc_hd__o211ai_1 _07598_ (.A1(_00040_),
    .A2(_00039_),
    .B1(_00052_),
    .C1(_00046_),
    .Y(_02689_));
 sky130_fd_sc_hd__a21oi_1 _07599_ (.A1(_02687_),
    .A2(_02688_),
    .B1(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__a21oi_1 _07600_ (.A1(_00062_),
    .A2(_00055_),
    .B1(_00061_),
    .Y(_02691_));
 sky130_fd_sc_hd__a21oi_1 _07601_ (.A1(_00052_),
    .A2(_00045_),
    .B1(_00051_),
    .Y(_02692_));
 sky130_fd_sc_hd__nand2_1 _07602_ (.A(_02691_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__nand2_1 _07603_ (.A(_00070_),
    .B(_00076_),
    .Y(_02694_));
 sky130_fd_sc_hd__a211oi_1 _07604_ (.A1(_02614_),
    .A2(_02691_),
    .B1(_02683_),
    .C1(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__o21ai_0 _07605_ (.A1(_02690_),
    .A2(_02693_),
    .B1(_02695_),
    .Y(_02696_));
 sky130_fd_sc_hd__nor2b_1 _07606_ (.A(_02686_),
    .B_N(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__xnor2_1 _07607_ (.A(_02682_),
    .B(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__nor4_1 _07608_ (.A(_00070_),
    .B(_00076_),
    .C(_00080_),
    .D(_00086_),
    .Y(_02699_));
 sky130_fd_sc_hd__nor2b_1 _07609_ (.A(_00034_),
    .B_N(_00007_),
    .Y(_02700_));
 sky130_fd_sc_hd__or2_2 _07610_ (.A(_00037_),
    .B(_00041_),
    .X(_02701_));
 sky130_fd_sc_hd__nand2b_1 _07611_ (.A_N(_00041_),
    .B(_00040_),
    .Y(_02702_));
 sky130_fd_sc_hd__nor2_1 _07612_ (.A(_00046_),
    .B(_00052_),
    .Y(_02703_));
 sky130_fd_sc_hd__o211ai_1 _07613_ (.A1(_02700_),
    .A2(_02701_),
    .B1(_02702_),
    .C1(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__nor2b_1 _07614_ (.A(_00052_),
    .B_N(_00047_),
    .Y(_02705_));
 sky130_fd_sc_hd__nor4_1 _07615_ (.A(_00053_),
    .B(_00057_),
    .C(_00063_),
    .D(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__inv_1 _07616_ (.A(_00062_),
    .Y(_02707_));
 sky130_fd_sc_hd__nand2b_1 _07617_ (.A_N(_00057_),
    .B(_00056_),
    .Y(_02708_));
 sky130_fd_sc_hd__a21oi_1 _07618_ (.A1(_02707_),
    .A2(_02708_),
    .B1(_00063_),
    .Y(_02709_));
 sky130_fd_sc_hd__a21oi_1 _07619_ (.A1(_02704_),
    .A2(_02706_),
    .B1(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__o21bai_1 _07620_ (.A1(_02601_),
    .A2(_00076_),
    .B1_N(_00077_),
    .Y(_02711_));
 sky130_fd_sc_hd__nor2b_1 _07621_ (.A(_00086_),
    .B_N(_00081_),
    .Y(_02712_));
 sky130_fd_sc_hd__a311o_1 _07622_ (.A1(_02592_),
    .A2(_02610_),
    .A3(_02711_),
    .B1(_02712_),
    .C1(_00087_),
    .X(_02713_));
 sky130_fd_sc_hd__a21oi_1 _07623_ (.A1(_02699_),
    .A2(_02710_),
    .B1(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__xnor2_1 _07624_ (.A(_00092_),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__a22oi_1 _07625_ (.A1(net477),
    .A2(_02698_),
    .B1(_02715_),
    .B2(net612),
    .Y(_02716_));
 sky130_fd_sc_hd__o2bb2ai_1 _07626_ (.A1_N(_02680_),
    .A2_N(_02716_),
    .B1(net557),
    .B2(_02666_),
    .Y(_02717_));
 sky130_fd_sc_hd__nor2_1 _07627_ (.A(net562),
    .B(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__or3_1 _07628_ (.A(\core.CPU_reset_a3 ),
    .B(_02650_),
    .C(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__nand3_1 _07630_ (.A(\core.CPU_Xreg_value_a4[10][11] ),
    .B(net550),
    .C(net428),
    .Y(_02721_));
 sky130_fd_sc_hd__o21ai_0 _07631_ (.A1(net428),
    .A2(net361),
    .B1(_02721_),
    .Y(_00754_));
 sky130_fd_sc_hd__a21o_1 _07634_ (.A1(_00092_),
    .A2(_00085_),
    .B1(_00091_),
    .X(_02724_));
 sky130_fd_sc_hd__a211oi_1 _07635_ (.A1(_02616_),
    .A2(_02623_),
    .B1(_02610_),
    .C1(_02682_),
    .Y(_02725_));
 sky130_fd_sc_hd__nor3_1 _07636_ (.A(_00098_),
    .B(_02724_),
    .C(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__o21ai_0 _07638_ (.A1(_02724_),
    .A2(_02725_),
    .B1(_00098_),
    .Y(_02728_));
 sky130_fd_sc_hd__nor3b_1 _07639_ (.A(_02726_),
    .B(net556),
    .C_N(_02728_),
    .Y(_02729_));
 sky130_fd_sc_hd__nand2_1 _07642_ (.A(_00089_),
    .B(_00095_),
    .Y(_02732_));
 sky130_fd_sc_hd__a21oi_1 _07643_ (.A1(_00083_),
    .A2(_00072_),
    .B1(_00082_),
    .Y(_02733_));
 sky130_fd_sc_hd__a21oi_1 _07644_ (.A1(_00095_),
    .A2(_00088_),
    .B1(_00094_),
    .Y(_02734_));
 sky130_fd_sc_hd__o21ai_0 _07645_ (.A1(_02732_),
    .A2(_02733_),
    .B1(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__nand4_1 _07646_ (.A(_00083_),
    .B(_00089_),
    .C(_00095_),
    .D(_00073_),
    .Y(_02736_));
 sky130_fd_sc_hd__a21oi_1 _07647_ (.A1(_02628_),
    .A2(_02634_),
    .B1(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__o21a_1 _07648_ (.A1(_02735_),
    .A2(_02737_),
    .B1(_00101_),
    .X(_02738_));
 sky130_fd_sc_hd__nor3_1 _07649_ (.A(_00101_),
    .B(_02735_),
    .C(_02737_),
    .Y(_02739_));
 sky130_fd_sc_hd__mux4_2 _07651_ (.A0(\core.CPU_src1_value_a3[5] ),
    .A1(\core.CPU_src1_value_a3[6] ),
    .A2(\core.CPU_src1_value_a3[7] ),
    .A3(\core.CPU_src1_value_a3[8] ),
    .S0(net554),
    .S1(net548),
    .X(_02741_));
 sky130_fd_sc_hd__mux4_2 _07653_ (.A0(\core.CPU_src1_value_a3[9] ),
    .A1(\core.CPU_src1_value_a3[10] ),
    .A2(\core.CPU_src1_value_a3[11] ),
    .A3(\core.CPU_src1_value_a3[12] ),
    .S0(net554),
    .S1(net548),
    .X(_02743_));
 sky130_fd_sc_hd__mux2i_1 _07655_ (.A0(_02741_),
    .A1(_02743_),
    .S(net553),
    .Y(_02745_));
 sky130_fd_sc_hd__mux4_2 _07657_ (.A0(\core.CPU_src1_value_a3[3] ),
    .A1(\core.CPU_src1_value_a3[1] ),
    .A2(\core.CPU_src1_value_a3[4] ),
    .A3(\core.CPU_src1_value_a3[2] ),
    .S0(_02577_),
    .S1(net554),
    .X(_02747_));
 sky130_fd_sc_hd__mux2i_1 _07658_ (.A0(net479),
    .A1(_02747_),
    .S(net553),
    .Y(_02748_));
 sky130_fd_sc_hd__mux2_2 _07660_ (.A0(_02745_),
    .A1(_02748_),
    .S(net480),
    .X(_02750_));
 sky130_fd_sc_hd__o32a_1 _07661_ (.A1(_02540_),
    .A2(_02738_),
    .A3(_02739_),
    .B1(_02750_),
    .B2(_02525_),
    .X(_02751_));
 sky130_fd_sc_hd__nor2_1 _07662_ (.A(net609),
    .B(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__a21oi_1 _07663_ (.A1(_02682_),
    .A2(_00087_),
    .B1(_00093_),
    .Y(_02753_));
 sky130_fd_sc_hd__inv_1 _07664_ (.A(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__or2_1 _07665_ (.A(_00086_),
    .B(_00092_),
    .X(_02755_));
 sky130_fd_sc_hd__a21oi_1 _07666_ (.A1(_02593_),
    .A2(_02606_),
    .B1(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__nor3_1 _07667_ (.A(_00098_),
    .B(_02754_),
    .C(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__o21ai_0 _07668_ (.A1(_02754_),
    .A2(_02756_),
    .B1(_00098_),
    .Y(_02758_));
 sky130_fd_sc_hd__nand3b_1 _07669_ (.A_N(_02757_),
    .B(net612),
    .C(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__o311ai_0 _07670_ (.A1(net612),
    .A2(_02729_),
    .A3(_02752_),
    .B1(_02759_),
    .C1(net557),
    .Y(_02760_));
 sky130_fd_sc_hd__nor2_1 _07673_ (.A(_02738_),
    .B(_02739_),
    .Y(_02763_));
 sky130_fd_sc_hd__a21oi_1 _07674_ (.A1(net611),
    .A2(_02763_),
    .B1(net562),
    .Y(_02764_));
 sky130_fd_sc_hd__nor2_1 _07676_ (.A(\core.CPU_dmem_rd_data_a5[12] ),
    .B(net536),
    .Y(_02766_));
 sky130_fd_sc_hd__a21oi_1 _07677_ (.A1(net370),
    .A2(_02764_),
    .B1(_02766_),
    .Y(_02767_));
 sky130_fd_sc_hd__nand2_1 _07678_ (.A(net429),
    .B(net360),
    .Y(_02768_));
 sky130_fd_sc_hd__nand2_1 _07679_ (.A(\core.CPU_Xreg_value_a4[10][12] ),
    .B(net428),
    .Y(_02769_));
 sky130_fd_sc_hd__a21oi_1 _07680_ (.A1(_02768_),
    .A2(_02769_),
    .B1(net607),
    .Y(_00755_));
 sky130_fd_sc_hd__nor2_1 _07681_ (.A(_02657_),
    .B(_02660_),
    .Y(_02770_));
 sky130_fd_sc_hd__o21ai_0 _07682_ (.A1(_02661_),
    .A2(_02770_),
    .B1(_02652_),
    .Y(_02771_));
 sky130_fd_sc_hd__a21oi_1 _07683_ (.A1(_00101_),
    .A2(_00094_),
    .B1(_00100_),
    .Y(_02772_));
 sky130_fd_sc_hd__nand2_1 _07684_ (.A(_02651_),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__nand2_1 _07685_ (.A(_00095_),
    .B(_00101_),
    .Y(_02774_));
 sky130_fd_sc_hd__a21oi_1 _07686_ (.A1(_02663_),
    .A2(_02662_),
    .B1(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__nand2b_1 _07687_ (.A_N(_02775_),
    .B(_02772_),
    .Y(_02776_));
 sky130_fd_sc_hd__o21ai_0 _07688_ (.A1(_02771_),
    .A2(_02773_),
    .B1(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__xnor2_1 _07689_ (.A(_00107_),
    .B(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__a21o_1 _07690_ (.A1(_00052_),
    .A2(_00045_),
    .B1(_00051_),
    .X(_02779_));
 sky130_fd_sc_hd__nor2_1 _07691_ (.A(_02694_),
    .B(_02614_),
    .Y(_02780_));
 sky130_fd_sc_hd__o21a_1 _07692_ (.A1(_02690_),
    .A2(_02779_),
    .B1(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__inv_1 _07693_ (.A(_00098_),
    .Y(_02782_));
 sky130_fd_sc_hd__a21oi_1 _07694_ (.A1(_00098_),
    .A2(_00091_),
    .B1(_00097_),
    .Y(_02783_));
 sky130_fd_sc_hd__o31ai_1 _07695_ (.A1(_02682_),
    .A2(_02782_),
    .A3(_02685_),
    .B1(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__o21ai_0 _07696_ (.A1(_02694_),
    .A2(_02691_),
    .B1(_02684_),
    .Y(_02785_));
 sky130_fd_sc_hd__or2_2 _07697_ (.A(_02784_),
    .B(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__nand4_1 _07698_ (.A(_00080_),
    .B(_00086_),
    .C(_00092_),
    .D(_00098_),
    .Y(_02787_));
 sky130_fd_sc_hd__nand2b_1 _07699_ (.A_N(_02784_),
    .B(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__o21ai_0 _07700_ (.A1(_02781_),
    .A2(_02786_),
    .B1(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__xnor2_1 _07701_ (.A(_00104_),
    .B(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__nor2_1 _07702_ (.A(net612),
    .B(net611),
    .Y(_02791_));
 sky130_fd_sc_hd__o21ai_0 _07703_ (.A1(net556),
    .A2(_02790_),
    .B1(net547),
    .Y(_02792_));
 sky130_fd_sc_hd__nand2_1 _07704_ (.A(net557),
    .B(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand2_1 _07705_ (.A(net557),
    .B(_02540_),
    .Y(_02794_));
 sky130_fd_sc_hd__mux4_2 _07706_ (.A0(\core.CPU_src1_value_a3[6] ),
    .A1(\core.CPU_src1_value_a3[7] ),
    .A2(\core.CPU_src1_value_a3[8] ),
    .A3(\core.CPU_src1_value_a3[9] ),
    .S0(net554),
    .S1(net548),
    .X(_02795_));
 sky130_fd_sc_hd__mux4_2 _07707_ (.A0(\core.CPU_src1_value_a3[10] ),
    .A1(\core.CPU_src1_value_a3[11] ),
    .A2(\core.CPU_src1_value_a3[12] ),
    .A3(\core.CPU_src1_value_a3[13] ),
    .S0(net554),
    .S1(net548),
    .X(_02796_));
 sky130_fd_sc_hd__mux2i_1 _07708_ (.A0(_02795_),
    .A1(_02796_),
    .S(net553),
    .Y(_02797_));
 sky130_fd_sc_hd__mux4_2 _07709_ (.A0(\core.CPU_src1_value_a3[2] ),
    .A1(\core.CPU_src1_value_a3[3] ),
    .A2(\core.CPU_src1_value_a3[4] ),
    .A3(\core.CPU_src1_value_a3[5] ),
    .S0(net554),
    .S1(net548),
    .X(_02798_));
 sky130_fd_sc_hd__mux2i_1 _07710_ (.A0(_00021_),
    .A1(_00003_),
    .S(_02570_),
    .Y(_02799_));
 sky130_fd_sc_hd__nand3_1 _07711_ (.A(net481),
    .B(net548),
    .C(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__a21boi_0 _07712_ (.A1(net553),
    .A2(_02798_),
    .B1_N(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__mux2_2 _07713_ (.A0(_02797_),
    .A1(_02801_),
    .S(net480),
    .X(_02802_));
 sky130_fd_sc_hd__o21a_1 _07714_ (.A1(_02525_),
    .A2(_02802_),
    .B1(net556),
    .X(_02803_));
 sky130_fd_sc_hd__nand2_1 _07715_ (.A(net612),
    .B(net557),
    .Y(_02804_));
 sky130_fd_sc_hd__a21oi_1 _07717_ (.A1(_02782_),
    .A2(_00093_),
    .B1(_00099_),
    .Y(_02806_));
 sky130_fd_sc_hd__o31ai_1 _07718_ (.A1(_00092_),
    .A2(_00098_),
    .A3(_02714_),
    .B1(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__xor2_1 _07719_ (.A(_00104_),
    .B(_02807_),
    .X(_02808_));
 sky130_fd_sc_hd__o22ai_1 _07720_ (.A1(_02792_),
    .A2(_02803_),
    .B1(_02804_),
    .B2(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__a31oi_1 _07721_ (.A1(_02778_),
    .A2(_02793_),
    .A3(_02794_),
    .B1(_02809_),
    .Y(_02810_));
 sky130_fd_sc_hd__and2_1 _07722_ (.A(net535),
    .B(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__o21ai_1 _07725_ (.A1(\core.CPU_dmem_rd_data_a5[13] ),
    .A2(net535),
    .B1(net551),
    .Y(_02814_));
 sky130_fd_sc_hd__nand3_1 _07729_ (.A(\core.CPU_Xreg_value_a4[10][13] ),
    .B(net552),
    .C(net428),
    .Y(_02818_));
 sky130_fd_sc_hd__o31ai_1 _07730_ (.A1(net428),
    .A2(_02811_),
    .A3(net439),
    .B1(_02818_),
    .Y(_00756_));
 sky130_fd_sc_hd__nor2_1 _07731_ (.A(net610),
    .B(\core.CPU_is_sll_a3 ),
    .Y(_02819_));
 sky130_fd_sc_hd__a221oi_1 _07732_ (.A1(_02629_),
    .A2(_02630_),
    .B1(_02631_),
    .B2(_02632_),
    .C1(_02633_),
    .Y(_02820_));
 sky130_fd_sc_hd__nand2_1 _07733_ (.A(_00101_),
    .B(_00107_),
    .Y(_02821_));
 sky130_fd_sc_hd__nor2_1 _07734_ (.A(_02736_),
    .B(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__nand2_1 _07735_ (.A(_02820_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _07736_ (.A(_00083_),
    .B(_00073_),
    .Y(_02824_));
 sky130_fd_sc_hd__o21ai_0 _07737_ (.A1(_02628_),
    .A2(_02824_),
    .B1(_02733_),
    .Y(_02825_));
 sky130_fd_sc_hd__nor2_1 _07738_ (.A(_02732_),
    .B(_02821_),
    .Y(_02826_));
 sky130_fd_sc_hd__a21oi_1 _07739_ (.A1(_00107_),
    .A2(_00100_),
    .B1(_00106_),
    .Y(_02827_));
 sky130_fd_sc_hd__o21ai_0 _07740_ (.A1(_02734_),
    .A2(_02821_),
    .B1(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__a21oi_1 _07741_ (.A1(_02825_),
    .A2(_02826_),
    .B1(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _07742_ (.A(_02823_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__xor2_1 _07743_ (.A(_00113_),
    .B(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_2 _07744_ (.A0(_02576_),
    .A1(_02575_),
    .S(net548),
    .X(_02832_));
 sky130_fd_sc_hd__mux4_2 _07745_ (.A0(\core.CPU_src1_value_a3[11] ),
    .A1(\core.CPU_src1_value_a3[12] ),
    .A2(\core.CPU_src1_value_a3[13] ),
    .A3(\core.CPU_src1_value_a3[14] ),
    .S0(net554),
    .S1(net548),
    .X(_02833_));
 sky130_fd_sc_hd__nand2_1 _07746_ (.A(net553),
    .B(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__o21ai_0 _07747_ (.A1(net553),
    .A2(_02832_),
    .B1(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__nand3_1 _07748_ (.A(net553),
    .B(_02577_),
    .C(_02573_),
    .Y(_02836_));
 sky130_fd_sc_hd__nand3_1 _07749_ (.A(net553),
    .B(_02572_),
    .C(net548),
    .Y(_02837_));
 sky130_fd_sc_hd__o211a_1 _07750_ (.A1(net553),
    .A2(_02586_),
    .B1(_02836_),
    .C1(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__mux2_2 _07751_ (.A0(_02835_),
    .A1(_02838_),
    .S(net480),
    .X(_02839_));
 sky130_fd_sc_hd__a221o_1 _07752_ (.A1(net546),
    .A2(_02831_),
    .B1(_02839_),
    .B2(_02667_),
    .C1(net609),
    .X(_02840_));
 sky130_fd_sc_hd__nor2_1 _07753_ (.A(_00056_),
    .B(_00055_),
    .Y(_02841_));
 sky130_fd_sc_hd__nor2_1 _07754_ (.A(_02707_),
    .B(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__o31a_1 _07755_ (.A1(_00051_),
    .A2(_00055_),
    .A3(_02613_),
    .B1(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__nand2_1 _07756_ (.A(_00098_),
    .B(_00104_),
    .Y(_02844_));
 sky130_fd_sc_hd__a21oi_1 _07757_ (.A1(_00092_),
    .A2(_00085_),
    .B1(_00091_),
    .Y(_02845_));
 sky130_fd_sc_hd__a21oi_1 _07758_ (.A1(_00104_),
    .A2(_00097_),
    .B1(_00103_),
    .Y(_02846_));
 sky130_fd_sc_hd__o21ai_0 _07759_ (.A1(_02844_),
    .A2(_02845_),
    .B1(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__o211ai_1 _07760_ (.A1(_02844_),
    .A2(_02845_),
    .B1(_02846_),
    .C1(_01146_),
    .Y(_02848_));
 sky130_fd_sc_hd__o211ai_1 _07761_ (.A1(_02844_),
    .A2(_02845_),
    .B1(_02846_),
    .C1(_01142_),
    .Y(_02849_));
 sky130_fd_sc_hd__o21a_1 _07762_ (.A1(_02622_),
    .A2(_02848_),
    .B1(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__o31a_1 _07763_ (.A1(_02622_),
    .A2(_02843_),
    .A3(_02847_),
    .B1(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__xnor2_1 _07764_ (.A(_00110_),
    .B(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hd__nand2_1 _07765_ (.A(net555),
    .B(net557),
    .Y(_02853_));
 sky130_fd_sc_hd__a21oi_1 _07766_ (.A1(net609),
    .A2(_02852_),
    .B1(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__inv_1 _07767_ (.A(_00110_),
    .Y(_02855_));
 sky130_fd_sc_hd__nand2b_1 _07768_ (.A_N(_00104_),
    .B(_00099_),
    .Y(_02856_));
 sky130_fd_sc_hd__nand2b_1 _07769_ (.A_N(_00105_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__or3_1 _07770_ (.A(_00098_),
    .B(_00104_),
    .C(_02755_),
    .X(_02858_));
 sky130_fd_sc_hd__o32ai_1 _07771_ (.A1(_00098_),
    .A2(_00104_),
    .A3(_02753_),
    .B1(_02858_),
    .B2(_02593_),
    .Y(_02859_));
 sky130_fd_sc_hd__nor3_1 _07772_ (.A(_00098_),
    .B(_00104_),
    .C(_02755_),
    .Y(_02860_));
 sky130_fd_sc_hd__o211a_1 _07773_ (.A1(_02598_),
    .A2(_02603_),
    .B1(_02860_),
    .C1(_02605_),
    .X(_02861_));
 sky130_fd_sc_hd__nor3_1 _07774_ (.A(_02857_),
    .B(net427),
    .C(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__xnor2_1 _07775_ (.A(_02855_),
    .B(_02862_),
    .Y(_02863_));
 sky130_fd_sc_hd__nor2_1 _07776_ (.A(net555),
    .B(net611),
    .Y(_02864_));
 sky130_fd_sc_hd__a22o_1 _07777_ (.A1(net611),
    .A2(_02831_),
    .B1(_02863_),
    .B2(net476),
    .X(_02865_));
 sky130_fd_sc_hd__a21oi_1 _07778_ (.A1(_02840_),
    .A2(_02854_),
    .B1(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__nand2_1 _07779_ (.A(net536),
    .B(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__o211ai_1 _07780_ (.A1(\core.CPU_dmem_rd_data_a5[14] ),
    .A2(net536),
    .B1(_02867_),
    .C1(_02644_),
    .Y(_02868_));
 sky130_fd_sc_hd__nand3_1 _07782_ (.A(\core.CPU_Xreg_value_a4[10][14] ),
    .B(net549),
    .C(net428),
    .Y(_02870_));
 sky130_fd_sc_hd__o21ai_0 _07783_ (.A1(net428),
    .A2(net347),
    .B1(_02870_),
    .Y(_00757_));
 sky130_fd_sc_hd__nand2_1 _07784_ (.A(_00104_),
    .B(_00110_),
    .Y(_02871_));
 sky130_fd_sc_hd__a21oi_1 _07785_ (.A1(_00110_),
    .A2(_00103_),
    .B1(_00109_),
    .Y(_02872_));
 sky130_fd_sc_hd__o21ai_0 _07786_ (.A1(_02783_),
    .A2(_02871_),
    .B1(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__nor2_1 _07787_ (.A(_02686_),
    .B(_02873_),
    .Y(_02874_));
 sky130_fd_sc_hd__nor3_1 _07788_ (.A(_00092_),
    .B(_00091_),
    .C(_00097_),
    .Y(_02875_));
 sky130_fd_sc_hd__nor2_1 _07789_ (.A(_00098_),
    .B(_00097_),
    .Y(_02876_));
 sky130_fd_sc_hd__o31ai_1 _07790_ (.A1(_02871_),
    .A2(_02875_),
    .A3(_02876_),
    .B1(_02872_),
    .Y(_02877_));
 sky130_fd_sc_hd__a21boi_0 _07791_ (.A1(_02696_),
    .A2(_02874_),
    .B1_N(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__xnor2_1 _07792_ (.A(_00116_),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__nand2_1 _07793_ (.A(_00107_),
    .B(_00113_),
    .Y(_02880_));
 sky130_fd_sc_hd__nand4_1 _07794_ (.A(_00095_),
    .B(_00101_),
    .C(_00107_),
    .D(_00113_),
    .Y(_02881_));
 sky130_fd_sc_hd__a21oi_1 _07795_ (.A1(_00113_),
    .A2(_00106_),
    .B1(_00112_),
    .Y(_02882_));
 sky130_fd_sc_hd__o211ai_1 _07796_ (.A1(_02772_),
    .A2(_02880_),
    .B1(_02881_),
    .C1(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__o21a_1 _07797_ (.A1(_02772_),
    .A2(_02880_),
    .B1(_02882_),
    .X(_02884_));
 sky130_fd_sc_hd__nand2_1 _07798_ (.A(net435),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__inv_1 _07799_ (.A(_00121_),
    .Y(_02886_));
 sky130_fd_sc_hd__a21oi_1 _07800_ (.A1(_02883_),
    .A2(_02885_),
    .B1(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__and3_1 _07801_ (.A(_02886_),
    .B(_02883_),
    .C(_02885_),
    .X(_02888_));
 sky130_fd_sc_hd__o21ai_0 _07802_ (.A1(_02887_),
    .A2(_02888_),
    .B1(net546),
    .Y(_02889_));
 sky130_fd_sc_hd__mux4_2 _07804_ (.A0(\core.CPU_src1_value_a3[12] ),
    .A1(\core.CPU_src1_value_a3[13] ),
    .A2(\core.CPU_src1_value_a3[14] ),
    .A3(\core.CPU_src1_value_a3[15] ),
    .S0(net554),
    .S1(net548),
    .X(_02891_));
 sky130_fd_sc_hd__mux2i_1 _07805_ (.A0(_02672_),
    .A1(_02891_),
    .S(net553),
    .Y(_02892_));
 sky130_fd_sc_hd__nand2_1 _07806_ (.A(net478),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__mux4_2 _07807_ (.A0(_02668_),
    .A1(_02669_),
    .A2(_02675_),
    .A3(_02676_),
    .S0(net554),
    .S1(net553),
    .X(_02894_));
 sky130_fd_sc_hd__nand2_1 _07808_ (.A(net480),
    .B(_02894_),
    .Y(_02895_));
 sky130_fd_sc_hd__a31oi_1 _07809_ (.A1(_02667_),
    .A2(_02893_),
    .A3(_02895_),
    .B1(net609),
    .Y(_02896_));
 sky130_fd_sc_hd__a221oi_1 _07810_ (.A1(net609),
    .A2(_02879_),
    .B1(_02889_),
    .B2(_02896_),
    .C1(_02853_),
    .Y(_02897_));
 sky130_fd_sc_hd__inv_1 _07811_ (.A(_00116_),
    .Y(_02898_));
 sky130_fd_sc_hd__nor4_1 _07812_ (.A(_00092_),
    .B(_00098_),
    .C(_00104_),
    .D(_00110_),
    .Y(_02899_));
 sky130_fd_sc_hd__nand2_1 _07813_ (.A(_02699_),
    .B(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__a211oi_1 _07814_ (.A1(_02704_),
    .A2(_02706_),
    .B1(_02709_),
    .C1(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__a21oi_1 _07815_ (.A1(_02855_),
    .A2(_00105_),
    .B1(_00111_),
    .Y(_02902_));
 sky130_fd_sc_hd__o31ai_1 _07816_ (.A1(_00104_),
    .A2(_00110_),
    .A3(_02806_),
    .B1(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__a21oi_1 _07817_ (.A1(_02713_),
    .A2(_02899_),
    .B1(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__nand2b_1 _07818_ (.A_N(_02901_),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__xnor2_1 _07819_ (.A(_02898_),
    .B(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__o21ai_0 _07820_ (.A1(_02887_),
    .A2(_02888_),
    .B1(net611),
    .Y(_02907_));
 sky130_fd_sc_hd__o21ai_0 _07821_ (.A1(_02804_),
    .A2(_02906_),
    .B1(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__nor2_1 _07822_ (.A(_02897_),
    .B(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__nor2_1 _07823_ (.A(\core.CPU_dmem_rd_data_a5[15] ),
    .B(net536),
    .Y(_02910_));
 sky130_fd_sc_hd__a211o_1 _07824_ (.A1(net535),
    .A2(_02909_),
    .B1(_02910_),
    .C1(\core.CPU_reset_a3 ),
    .X(_02911_));
 sky130_fd_sc_hd__nand3_1 _07827_ (.A(\core.CPU_Xreg_value_a4[10][15] ),
    .B(net551),
    .C(_02563_),
    .Y(_02914_));
 sky130_fd_sc_hd__o21ai_0 _07828_ (.A1(_02563_),
    .A2(_02911_),
    .B1(_02914_),
    .Y(_00758_));
 sky130_fd_sc_hd__nor2_1 _07829_ (.A(net609),
    .B(_02540_),
    .Y(_02915_));
 sky130_fd_sc_hd__inv_1 _07830_ (.A(\core.CPU_imm_a3[5] ),
    .Y(_02916_));
 sky130_fd_sc_hd__mux2i_1 _07831_ (.A0(\core.CPU_is_sll_a3 ),
    .A1(_02916_),
    .S(net610),
    .Y(_02917_));
 sky130_fd_sc_hd__nand2_1 _07832_ (.A(net610),
    .B(\core.CPU_imm_a3[4] ),
    .Y(_02918_));
 sky130_fd_sc_hd__o21ai_0 _07833_ (.A1(net610),
    .A2(_00050_),
    .B1(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__nor3_1 _07834_ (.A(net609),
    .B(net475),
    .C(net474),
    .Y(_02920_));
 sky130_fd_sc_hd__mux2i_1 _07835_ (.A0(_02741_),
    .A1(_02747_),
    .S(net481),
    .Y(_02921_));
 sky130_fd_sc_hd__nand2_1 _07836_ (.A(net480),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__nand2_1 _07837_ (.A(net481),
    .B(_02743_),
    .Y(_02923_));
 sky130_fd_sc_hd__mux4_2 _07839_ (.A0(\core.CPU_src1_value_a3[13] ),
    .A1(\core.CPU_src1_value_a3[14] ),
    .A2(\core.CPU_src1_value_a3[15] ),
    .A3(\core.CPU_src1_value_a3[16] ),
    .S0(net554),
    .S1(net548),
    .X(_02925_));
 sky130_fd_sc_hd__nand2_1 _07840_ (.A(net553),
    .B(_02925_),
    .Y(_02926_));
 sky130_fd_sc_hd__nand3_1 _07841_ (.A(net478),
    .B(_02923_),
    .C(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__nand3_1 _07842_ (.A(_02920_),
    .B(_02922_),
    .C(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__nor2_1 _07843_ (.A(net609),
    .B(net475),
    .Y(_02929_));
 sky130_fd_sc_hd__nand3b_1 _07844_ (.A_N(\core.CPU_imm_a3[3] ),
    .B(\core.CPU_imm_a3[4] ),
    .C(net610),
    .Y(_02930_));
 sky130_fd_sc_hd__o41ai_1 _07845_ (.A1(net610),
    .A2(\core.CPU_src2_value_a3[2] ),
    .A3(\core.CPU_src2_value_a3[3] ),
    .A4(_00050_),
    .B1(_02930_),
    .Y(_02931_));
 sky130_fd_sc_hd__nand3_1 _07846_ (.A(net479),
    .B(_02929_),
    .C(net473),
    .Y(_02932_));
 sky130_fd_sc_hd__nand3_1 _07847_ (.A(net547),
    .B(_02928_),
    .C(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2b_1 _07848_ (.A_N(_00124_),
    .B(net609),
    .Y(_02934_));
 sky130_fd_sc_hd__nand2_1 _07849_ (.A(net609),
    .B(_00124_),
    .Y(_02935_));
 sky130_fd_sc_hd__nor3_1 _07850_ (.A(_02855_),
    .B(_02898_),
    .C(_01142_),
    .Y(_02936_));
 sky130_fd_sc_hd__a21oi_1 _07851_ (.A1(_00110_),
    .A2(_02847_),
    .B1(_00109_),
    .Y(_02937_));
 sky130_fd_sc_hd__nor2_1 _07852_ (.A(_02898_),
    .B(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__a211oi_1 _07853_ (.A1(_02624_),
    .A2(_02936_),
    .B1(_02938_),
    .C1(_00115_),
    .Y(_02939_));
 sky130_fd_sc_hd__mux2i_1 _07854_ (.A0(_02934_),
    .A1(_02935_),
    .S(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__a21oi_1 _07855_ (.A1(_00121_),
    .A2(_00112_),
    .B1(_00120_),
    .Y(_02941_));
 sky130_fd_sc_hd__nand2_1 _07856_ (.A(_00113_),
    .B(_00121_),
    .Y(_02942_));
 sky130_fd_sc_hd__a21o_1 _07857_ (.A1(_02823_),
    .A2(_02829_),
    .B1(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__nand2_1 _07858_ (.A(_02941_),
    .B(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__xor2_1 _07859_ (.A(_00119_),
    .B(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__o31ai_1 _07860_ (.A1(_02915_),
    .A2(_02933_),
    .A3(_02940_),
    .B1(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__o21ai_0 _07861_ (.A1(_02933_),
    .A2(_02940_),
    .B1(net557),
    .Y(_02947_));
 sky130_fd_sc_hd__nor2_1 _07862_ (.A(net427),
    .B(_02861_),
    .Y(_02948_));
 sky130_fd_sc_hd__inv_1 _07863_ (.A(_00111_),
    .Y(_02949_));
 sky130_fd_sc_hd__nor2_1 _07864_ (.A(_00105_),
    .B(_00111_),
    .Y(_02950_));
 sky130_fd_sc_hd__a221oi_1 _07865_ (.A1(_00110_),
    .A2(_02949_),
    .B1(_02856_),
    .B2(_02950_),
    .C1(_00116_),
    .Y(_02951_));
 sky130_fd_sc_hd__nor2_1 _07866_ (.A(_00117_),
    .B(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__o31ai_1 _07867_ (.A1(_00110_),
    .A2(_00116_),
    .A3(_02948_),
    .B1(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__xor2_1 _07868_ (.A(_00124_),
    .B(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__a22oi_1 _07870_ (.A1(_02946_),
    .A2(_02947_),
    .B1(_02954_),
    .B2(net476),
    .Y(_02956_));
 sky130_fd_sc_hd__mux2i_1 _07871_ (.A0(\core.CPU_dmem_rd_data_a5[16] ),
    .A1(_02956_),
    .S(net535),
    .Y(_02957_));
 sky130_fd_sc_hd__o21ai_0 _07874_ (.A1(\core.CPU_Xreg_value_a4[10][16] ),
    .A2(net429),
    .B1(net551),
    .Y(_02960_));
 sky130_fd_sc_hd__a21oi_1 _07875_ (.A1(net429),
    .A2(net346),
    .B1(_02960_),
    .Y(_00759_));
 sky130_fd_sc_hd__nor2_1 _07876_ (.A(\core.CPU_reset_a3 ),
    .B(_01114_),
    .Y(_02961_));
 sky130_fd_sc_hd__nand2_1 _07877_ (.A(net429),
    .B(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__o21bai_1 _07878_ (.A1(_02886_),
    .A2(_02882_),
    .B1_N(_00120_),
    .Y(_02963_));
 sky130_fd_sc_hd__a21oi_1 _07879_ (.A1(_00119_),
    .A2(_02963_),
    .B1(_00118_),
    .Y(_02964_));
 sky130_fd_sc_hd__o21ai_0 _07880_ (.A1(_02651_),
    .A2(_02774_),
    .B1(_02772_),
    .Y(_02965_));
 sky130_fd_sc_hd__nand2_1 _07881_ (.A(_00121_),
    .B(_00119_),
    .Y(_02966_));
 sky130_fd_sc_hd__nor2_1 _07882_ (.A(_02880_),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__o211ai_1 _07883_ (.A1(_02771_),
    .A2(_02965_),
    .B1(_02967_),
    .C1(_02776_),
    .Y(_02968_));
 sky130_fd_sc_hd__nand2_1 _07884_ (.A(_02964_),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__xnor2_1 _07885_ (.A(_00127_),
    .B(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__inv_1 _07887_ (.A(_00130_),
    .Y(_02972_));
 sky130_fd_sc_hd__a21oi_1 _07888_ (.A1(_00124_),
    .A2(_00115_),
    .B1(_00123_),
    .Y(_02973_));
 sky130_fd_sc_hd__inv_1 _07889_ (.A(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__a31oi_1 _07890_ (.A1(_00116_),
    .A2(_00124_),
    .A3(_02878_),
    .B1(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__xnor2_1 _07891_ (.A(_02972_),
    .B(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__nand2_1 _07892_ (.A(net609),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__a31oi_1 _07893_ (.A1(net555),
    .A2(net546),
    .A3(_02977_),
    .B1(net611),
    .Y(_02978_));
 sky130_fd_sc_hd__nand2_1 _07894_ (.A(net556),
    .B(_02791_),
    .Y(_02979_));
 sky130_fd_sc_hd__nor2b_1 _07896_ (.A(net610),
    .B_N(\core.CPU_src2_value_a3[4] ),
    .Y(_02981_));
 sky130_fd_sc_hd__a21oi_1 _07897_ (.A1(net610),
    .A2(\core.CPU_imm_a3[4] ),
    .B1(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__mux4_2 _07898_ (.A0(\core.CPU_src1_value_a3[14] ),
    .A1(\core.CPU_src1_value_a3[15] ),
    .A2(\core.CPU_src1_value_a3[16] ),
    .A3(\core.CPU_src1_value_a3[17] ),
    .S0(net554),
    .S1(net548),
    .X(_02983_));
 sky130_fd_sc_hd__nand2_1 _07899_ (.A(_02982_),
    .B(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__a31oi_1 _07901_ (.A1(net474),
    .A2(net548),
    .A3(_02799_),
    .B1(net481),
    .Y(_02986_));
 sky130_fd_sc_hd__a21oi_1 _07902_ (.A1(_02982_),
    .A2(_02796_),
    .B1(net553),
    .Y(_02987_));
 sky130_fd_sc_hd__a21oi_1 _07903_ (.A1(_02984_),
    .A2(_02986_),
    .B1(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__mux2i_1 _07904_ (.A0(_02795_),
    .A1(_02798_),
    .S(net481),
    .Y(_02989_));
 sky130_fd_sc_hd__nand2_1 _07905_ (.A(_02982_),
    .B(net480),
    .Y(_02990_));
 sky130_fd_sc_hd__nor2_1 _07906_ (.A(_02989_),
    .B(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__a21oi_1 _07907_ (.A1(net478),
    .A2(_02988_),
    .B1(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__o31ai_1 _07908_ (.A1(net475),
    .A2(_02979_),
    .A3(_02992_),
    .B1(_02976_),
    .Y(_02993_));
 sky130_fd_sc_hd__nand2_1 _07909_ (.A(net609),
    .B(net547),
    .Y(_02994_));
 sky130_fd_sc_hd__o31ai_1 _07910_ (.A1(net475),
    .A2(_02853_),
    .A3(_02992_),
    .B1(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__nor4_1 _07911_ (.A(_00104_),
    .B(_00110_),
    .C(_00116_),
    .D(_00124_),
    .Y(_02996_));
 sky130_fd_sc_hd__nor2b_1 _07912_ (.A(_00124_),
    .B_N(_00117_),
    .Y(_02997_));
 sky130_fd_sc_hd__nor2_1 _07913_ (.A(_00125_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__o31ai_1 _07914_ (.A1(_00116_),
    .A2(_00124_),
    .A3(_02902_),
    .B1(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__a21oi_1 _07915_ (.A1(_02807_),
    .A2(_02996_),
    .B1(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__xnor2_1 _07916_ (.A(_02972_),
    .B(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__a22oi_1 _07917_ (.A1(_02993_),
    .A2(_02995_),
    .B1(_03001_),
    .B2(net476),
    .Y(_03002_));
 sky130_fd_sc_hd__o21a_1 _07918_ (.A1(_02970_),
    .A2(_02978_),
    .B1(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__nand3_1 _07921_ (.A(net551),
    .B(\core.CPU_dmem_rd_data_a5[17] ),
    .C(_01114_),
    .Y(_03006_));
 sky130_fd_sc_hd__nor2_1 _07923_ (.A(net428),
    .B(_03006_),
    .Y(_03008_));
 sky130_fd_sc_hd__a31oi_1 _07924_ (.A1(\core.CPU_Xreg_value_a4[10][17] ),
    .A2(net552),
    .A3(net428),
    .B1(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__o21ai_0 _07925_ (.A1(_02962_),
    .A2(_03003_),
    .B1(_03009_),
    .Y(_00760_));
 sky130_fd_sc_hd__mux4_2 _07926_ (.A0(\core.CPU_src1_value_a3[15] ),
    .A1(\core.CPU_src1_value_a3[16] ),
    .A2(\core.CPU_src1_value_a3[17] ),
    .A3(\core.CPU_src1_value_a3[18] ),
    .S0(net554),
    .S1(net548),
    .X(_03010_));
 sky130_fd_sc_hd__mux2i_1 _07927_ (.A0(_02833_),
    .A1(_03010_),
    .S(net553),
    .Y(_03011_));
 sky130_fd_sc_hd__mux2i_1 _07928_ (.A0(_02580_),
    .A1(_03011_),
    .S(net478),
    .Y(_03012_));
 sky130_fd_sc_hd__a221oi_1 _07929_ (.A1(_02586_),
    .A2(net473),
    .B1(_03012_),
    .B2(_02982_),
    .C1(net546),
    .Y(_03013_));
 sky130_fd_sc_hd__inv_1 _07930_ (.A(_00133_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand2_1 _07931_ (.A(_00119_),
    .B(_00127_),
    .Y(_03015_));
 sky130_fd_sc_hd__a21oi_1 _07932_ (.A1(_00127_),
    .A2(_00118_),
    .B1(_00126_),
    .Y(_03016_));
 sky130_fd_sc_hd__o21ai_0 _07933_ (.A1(_02941_),
    .A2(_03015_),
    .B1(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hd__nand4_1 _07934_ (.A(_00113_),
    .B(_00121_),
    .C(_00119_),
    .D(_00127_),
    .Y(_03018_));
 sky130_fd_sc_hd__a21oi_1 _07935_ (.A1(_02823_),
    .A2(_02829_),
    .B1(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__nor2_1 _07936_ (.A(_03017_),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__xnor2_1 _07937_ (.A(_03014_),
    .B(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__o22ai_1 _07938_ (.A1(net475),
    .A2(_03013_),
    .B1(_03021_),
    .B2(_02540_),
    .Y(_03022_));
 sky130_fd_sc_hd__nand2_1 _07939_ (.A(_00116_),
    .B(_00124_),
    .Y(_03023_));
 sky130_fd_sc_hd__nor3_1 _07940_ (.A(_02855_),
    .B(_02972_),
    .C(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__a211oi_1 _07941_ (.A1(_00116_),
    .A2(_00109_),
    .B1(_00115_),
    .C1(_00123_),
    .Y(_03025_));
 sky130_fd_sc_hd__o21ai_0 _07942_ (.A1(_00124_),
    .A2(_00123_),
    .B1(_00130_),
    .Y(_03026_));
 sky130_fd_sc_hd__inv_1 _07943_ (.A(_00129_),
    .Y(_03027_));
 sky130_fd_sc_hd__o21ai_0 _07944_ (.A1(_03025_),
    .A2(_03026_),
    .B1(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__a21oi_1 _07945_ (.A1(_03024_),
    .A2(_02851_),
    .B1(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__xor2_1 _07946_ (.A(_00136_),
    .B(_03029_),
    .X(_03030_));
 sky130_fd_sc_hd__a21oi_1 _07947_ (.A1(net609),
    .A2(_03030_),
    .B1(_02853_),
    .Y(_03031_));
 sky130_fd_sc_hd__or2_2 _07948_ (.A(_00124_),
    .B(_00130_),
    .X(_03032_));
 sky130_fd_sc_hd__a21oi_1 _07949_ (.A1(_02898_),
    .A2(_00111_),
    .B1(_00117_),
    .Y(_03033_));
 sky130_fd_sc_hd__nor3_1 _07950_ (.A(_00110_),
    .B(_00116_),
    .C(_03032_),
    .Y(_03034_));
 sky130_fd_sc_hd__o31ai_1 _07951_ (.A1(_02857_),
    .A2(net427),
    .A3(_02861_),
    .B1(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__nor2b_1 _07952_ (.A(_00130_),
    .B_N(_00125_),
    .Y(_03036_));
 sky130_fd_sc_hd__nor2_1 _07953_ (.A(_00131_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__o211ai_1 _07954_ (.A1(_03032_),
    .A2(_03033_),
    .B1(_03035_),
    .C1(_03037_),
    .Y(_03038_));
 sky130_fd_sc_hd__xnor2_1 _07955_ (.A(_00136_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__a2bb2oi_1 _07956_ (.A1_N(net557),
    .A2_N(_03021_),
    .B1(_03039_),
    .B2(net476),
    .Y(_03040_));
 sky130_fd_sc_hd__o21ai_0 _07957_ (.A1(_02994_),
    .A2(_03030_),
    .B1(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__a21oi_1 _07958_ (.A1(_03022_),
    .A2(_03031_),
    .B1(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__nand3_1 _07959_ (.A(net551),
    .B(\core.CPU_dmem_rd_data_a5[18] ),
    .C(_01114_),
    .Y(_03043_));
 sky130_fd_sc_hd__nand3_1 _07962_ (.A(\core.CPU_Xreg_value_a4[10][18] ),
    .B(net552),
    .C(net428),
    .Y(_03046_));
 sky130_fd_sc_hd__o221ai_1 _07963_ (.A1(_02962_),
    .A2(net359),
    .B1(_03043_),
    .B2(net428),
    .C1(_03046_),
    .Y(_00761_));
 sky130_fd_sc_hd__nor4_1 _07965_ (.A(_00116_),
    .B(_00124_),
    .C(_00130_),
    .D(_00136_),
    .Y(_03048_));
 sky130_fd_sc_hd__nor2_1 _07966_ (.A(_00130_),
    .B(_00136_),
    .Y(_03049_));
 sky130_fd_sc_hd__o21ai_0 _07967_ (.A1(_00125_),
    .A2(_02997_),
    .B1(_03049_),
    .Y(_03050_));
 sky130_fd_sc_hd__nor2b_1 _07968_ (.A(_00136_),
    .B_N(_00131_),
    .Y(_03051_));
 sky130_fd_sc_hd__nor2_1 _07969_ (.A(_00137_),
    .B(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__nand2_1 _07970_ (.A(_03050_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__a21oi_1 _07971_ (.A1(_02905_),
    .A2(net438),
    .B1(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__xnor2_1 _07972_ (.A(_00142_),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__inv_1 _07973_ (.A(_00142_),
    .Y(_03056_));
 sky130_fd_sc_hd__nand2_1 _07974_ (.A(_00130_),
    .B(_00136_),
    .Y(_03057_));
 sky130_fd_sc_hd__o21a_1 _07975_ (.A1(_03023_),
    .A2(_02872_),
    .B1(_02973_),
    .X(_03058_));
 sky130_fd_sc_hd__a21oi_1 _07976_ (.A1(_00136_),
    .A2(_00129_),
    .B1(_00135_),
    .Y(_03059_));
 sky130_fd_sc_hd__o21a_1 _07977_ (.A1(_03057_),
    .A2(_03058_),
    .B1(_03059_),
    .X(_03060_));
 sky130_fd_sc_hd__inv_1 _07978_ (.A(_02871_),
    .Y(_03061_));
 sky130_fd_sc_hd__nor2_1 _07979_ (.A(_03023_),
    .B(_03057_),
    .Y(_03062_));
 sky130_fd_sc_hd__o2111ai_1 _07980_ (.A1(_02781_),
    .A2(_02786_),
    .B1(_03061_),
    .C1(_03062_),
    .D1(_02788_),
    .Y(_03063_));
 sky130_fd_sc_hd__and3_1 _07981_ (.A(_03056_),
    .B(_03060_),
    .C(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__a21oi_1 _07982_ (.A1(_03060_),
    .A2(_03063_),
    .B1(_03056_),
    .Y(_03065_));
 sky130_fd_sc_hd__nand2_1 _07983_ (.A(net478),
    .B(_02891_),
    .Y(_03066_));
 sky130_fd_sc_hd__o211ai_1 _07984_ (.A1(net478),
    .A2(_02677_),
    .B1(_03066_),
    .C1(net481),
    .Y(_03067_));
 sky130_fd_sc_hd__mux4_2 _07985_ (.A0(\core.CPU_src1_value_a3[16] ),
    .A1(\core.CPU_src1_value_a3[17] ),
    .A2(\core.CPU_src1_value_a3[18] ),
    .A3(\core.CPU_src1_value_a3[19] ),
    .S0(net554),
    .S1(net548),
    .X(_03068_));
 sky130_fd_sc_hd__nand2_1 _07986_ (.A(net478),
    .B(_03068_),
    .Y(_03069_));
 sky130_fd_sc_hd__nand2_1 _07987_ (.A(net480),
    .B(_02672_),
    .Y(_03070_));
 sky130_fd_sc_hd__nand3_1 _07988_ (.A(net553),
    .B(_03069_),
    .C(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__a31o_2 _07989_ (.A1(_02670_),
    .A2(_02929_),
    .A3(net473),
    .B1(_02853_),
    .X(_03072_));
 sky130_fd_sc_hd__a31oi_1 _07990_ (.A1(_02920_),
    .A2(_03067_),
    .A3(_03071_),
    .B1(_03072_),
    .Y(_03073_));
 sky130_fd_sc_hd__o31ai_1 _07991_ (.A1(net556),
    .A2(_03064_),
    .A3(_03065_),
    .B1(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _07993_ (.A(_00127_),
    .B(_00133_),
    .Y(_03076_));
 sky130_fd_sc_hd__nor2_1 _07994_ (.A(_02966_),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__nand2_1 _07995_ (.A(_02883_),
    .B(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__o21ai_0 _07996_ (.A1(_02772_),
    .A2(_02880_),
    .B1(_02882_),
    .Y(_03079_));
 sky130_fd_sc_hd__a21oi_1 _07997_ (.A1(_00119_),
    .A2(_00120_),
    .B1(_00118_),
    .Y(_03080_));
 sky130_fd_sc_hd__a21oi_1 _07998_ (.A1(_00133_),
    .A2(_00126_),
    .B1(_00132_),
    .Y(_03081_));
 sky130_fd_sc_hd__o21ai_0 _07999_ (.A1(_03080_),
    .A2(_03076_),
    .B1(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__a21oi_1 _08000_ (.A1(_03079_),
    .A2(_03077_),
    .B1(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__o21ai_0 _08001_ (.A1(net435),
    .A2(_03078_),
    .B1(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__xnor2_1 _08002_ (.A(_00139_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_1 _08003_ (.A(net611),
    .B(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__nand2_1 _08004_ (.A(net556),
    .B(net546),
    .Y(_03087_));
 sky130_fd_sc_hd__nor2_1 _08005_ (.A(_03087_),
    .B(_03085_),
    .Y(_03088_));
 sky130_fd_sc_hd__a21oi_1 _08006_ (.A1(net376),
    .A2(_03086_),
    .B1(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__a211oi_1 _08007_ (.A1(net476),
    .A2(_03055_),
    .B1(_03089_),
    .C1(net562),
    .Y(_03090_));
 sky130_fd_sc_hd__a21oi_1 _08008_ (.A1(\core.CPU_dmem_rd_data_a5[19] ),
    .A2(net562),
    .B1(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__o21ai_0 _08009_ (.A1(\core.CPU_Xreg_value_a4[10][19] ),
    .A2(net429),
    .B1(_02644_),
    .Y(_03092_));
 sky130_fd_sc_hd__a21oi_1 _08010_ (.A1(net429),
    .A2(net358),
    .B1(_03092_),
    .Y(_00762_));
 sky130_fd_sc_hd__a32o_1 _08012_ (.A1(_02530_),
    .A2(net548),
    .A3(_02799_),
    .B1(net546),
    .B2(_00002_),
    .X(_03094_));
 sky130_fd_sc_hd__nand2_1 _08013_ (.A(net609),
    .B(_00006_),
    .Y(_03095_));
 sky130_fd_sc_hd__o21ai_0 _08014_ (.A1(net609),
    .A2(_03094_),
    .B1(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__nand2_1 _08015_ (.A(net612),
    .B(_00009_),
    .Y(_03097_));
 sky130_fd_sc_hd__o21ai_0 _08016_ (.A1(net612),
    .A2(_03096_),
    .B1(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__mux2_2 _08017_ (.A0(_00002_),
    .A1(_03098_),
    .S(net557),
    .X(_03099_));
 sky130_fd_sc_hd__mux2i_2 _08018_ (.A0(\core.CPU_dmem_rd_data_a5[1] ),
    .A1(_03099_),
    .S(net536),
    .Y(_03100_));
 sky130_fd_sc_hd__nor3_1 _08019_ (.A(\core.CPU_Xreg_value_a4[10][1] ),
    .B(net607),
    .C(_02558_),
    .Y(_03101_));
 sky130_fd_sc_hd__a31oi_1 _08020_ (.A1(_02644_),
    .A2(_02558_),
    .A3(net375),
    .B1(_03101_),
    .Y(_00763_));
 sky130_fd_sc_hd__mux4_2 _08021_ (.A0(\core.CPU_src1_value_a3[17] ),
    .A1(\core.CPU_src1_value_a3[18] ),
    .A2(\core.CPU_src1_value_a3[19] ),
    .A3(\core.CPU_src1_value_a3[20] ),
    .S0(net554),
    .S1(net548),
    .X(_03102_));
 sky130_fd_sc_hd__mux2i_1 _08022_ (.A0(_02925_),
    .A1(_03102_),
    .S(net553),
    .Y(_03103_));
 sky130_fd_sc_hd__nand2_1 _08023_ (.A(_02982_),
    .B(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__nand2_1 _08024_ (.A(net474),
    .B(_02748_),
    .Y(_03105_));
 sky130_fd_sc_hd__nor2_1 _08025_ (.A(_02745_),
    .B(_02990_),
    .Y(_03106_));
 sky130_fd_sc_hd__a31oi_1 _08026_ (.A1(net478),
    .A2(_03104_),
    .A3(_03105_),
    .B1(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__nor4_1 _08027_ (.A(_01127_),
    .B(_01130_),
    .C(_01142_),
    .D(_01146_),
    .Y(_03108_));
 sky130_fd_sc_hd__o311ai_0 _08028_ (.A1(_00051_),
    .A2(_00055_),
    .A3(_02613_),
    .B1(_02842_),
    .C1(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__nor2_1 _08029_ (.A(_01127_),
    .B(_02846_),
    .Y(_03110_));
 sky130_fd_sc_hd__a21oi_1 _08030_ (.A1(_00142_),
    .A2(_00135_),
    .B1(_00141_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand2_1 _08031_ (.A(_01130_),
    .B(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__o41ai_1 _08032_ (.A1(_00135_),
    .A2(_00141_),
    .A3(_03028_),
    .A4(_03110_),
    .B1(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__nor3_1 _08033_ (.A(_01127_),
    .B(_01130_),
    .C(_01142_),
    .Y(_03114_));
 sky130_fd_sc_hd__nor4_1 _08034_ (.A(_01127_),
    .B(_01130_),
    .C(_02844_),
    .D(_02845_),
    .Y(_03115_));
 sky130_fd_sc_hd__a21oi_1 _08035_ (.A1(_02622_),
    .A2(_03114_),
    .B1(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__nand3_1 _08036_ (.A(net393),
    .B(_03113_),
    .C(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__a211o_1 _08037_ (.A1(_03037_),
    .A2(_03032_),
    .B1(_00136_),
    .C1(_00142_),
    .X(_03118_));
 sky130_fd_sc_hd__nor4_1 _08038_ (.A(_00117_),
    .B(_00131_),
    .C(_02951_),
    .D(_03036_),
    .Y(_03119_));
 sky130_fd_sc_hd__nor2b_1 _08039_ (.A(_00142_),
    .B_N(_00137_),
    .Y(_03120_));
 sky130_fd_sc_hd__nor2_1 _08040_ (.A(_00143_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__o21a_1 _08041_ (.A1(_03118_),
    .A2(_03119_),
    .B1(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__nor2_1 _08042_ (.A(_00136_),
    .B(_00142_),
    .Y(_03123_));
 sky130_fd_sc_hd__o211ai_1 _08043_ (.A1(net427),
    .A2(_02861_),
    .B1(_03034_),
    .C1(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__and2_1 _08044_ (.A(_03122_),
    .B(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__o221ai_1 _08045_ (.A1(_02994_),
    .A2(_03117_),
    .B1(_03125_),
    .B2(_02804_),
    .C1(_00148_),
    .Y(_03126_));
 sky130_fd_sc_hd__nor2_1 _08046_ (.A(net611),
    .B(_02609_),
    .Y(_03127_));
 sky130_fd_sc_hd__a221o_1 _08047_ (.A1(_03127_),
    .A2(_03117_),
    .B1(_03125_),
    .B2(net476),
    .C1(_00148_),
    .X(_03128_));
 sky130_fd_sc_hd__o21ai_0 _08048_ (.A1(_02827_),
    .A2(_02942_),
    .B1(_02941_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_1 _08049_ (.A(_00133_),
    .B(_00139_),
    .Y(_03130_));
 sky130_fd_sc_hd__nor2_1 _08050_ (.A(_03015_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__inv_1 _08051_ (.A(_00139_),
    .Y(_03132_));
 sky130_fd_sc_hd__a21oi_1 _08052_ (.A1(_00139_),
    .A2(_00132_),
    .B1(_00138_),
    .Y(_03133_));
 sky130_fd_sc_hd__o31ai_1 _08053_ (.A1(_03014_),
    .A2(_03132_),
    .A3(_03016_),
    .B1(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__a21o_1 _08054_ (.A1(_03129_),
    .A2(_03131_),
    .B1(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__nor3_1 _08055_ (.A(_02821_),
    .B(_03018_),
    .C(_03130_),
    .Y(_03136_));
 sky130_fd_sc_hd__o21a_1 _08056_ (.A1(_02735_),
    .A2(_02737_),
    .B1(_03136_),
    .X(_03137_));
 sky130_fd_sc_hd__nor2_1 _08057_ (.A(_03135_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__xnor2_1 _08058_ (.A(_00145_),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__a22oi_1 _08059_ (.A1(_03126_),
    .A2(_03128_),
    .B1(_03139_),
    .B2(_02542_),
    .Y(_03140_));
 sky130_fd_sc_hd__o31ai_1 _08060_ (.A1(net475),
    .A2(_02979_),
    .A3(_03107_),
    .B1(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand2b_1 _08061_ (.A_N(\core.CPU_dmem_rd_data_a5[20] ),
    .B(net562),
    .Y(_03142_));
 sky130_fd_sc_hd__o211ai_1 _08062_ (.A1(net562),
    .A2(_03141_),
    .B1(_03142_),
    .C1(_02644_),
    .Y(_03143_));
 sky130_fd_sc_hd__nand3_1 _08064_ (.A(\core.CPU_Xreg_value_a4[10][20] ),
    .B(net549),
    .C(net428),
    .Y(_03145_));
 sky130_fd_sc_hd__o21ai_0 _08065_ (.A1(net428),
    .A2(net357),
    .B1(_03145_),
    .Y(_00764_));
 sky130_fd_sc_hd__inv_1 _08066_ (.A(_00154_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand4_1 _08067_ (.A(_00116_),
    .B(_00124_),
    .C(_00130_),
    .D(_00136_),
    .Y(_03147_));
 sky130_fd_sc_hd__nand2_1 _08068_ (.A(_00142_),
    .B(_00148_),
    .Y(_03148_));
 sky130_fd_sc_hd__nor4_1 _08069_ (.A(_02787_),
    .B(_02871_),
    .C(_03147_),
    .D(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__nor3_1 _08070_ (.A(_02871_),
    .B(_03147_),
    .C(_03148_),
    .Y(_03150_));
 sky130_fd_sc_hd__a22o_1 _08071_ (.A1(_02784_),
    .A2(_03150_),
    .B1(_03149_),
    .B2(_02785_),
    .X(_03151_));
 sky130_fd_sc_hd__a21o_1 _08072_ (.A1(_02781_),
    .A2(_03149_),
    .B1(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__a21oi_1 _08073_ (.A1(_00148_),
    .A2(_00141_),
    .B1(_00147_),
    .Y(_03153_));
 sky130_fd_sc_hd__o21a_1 _08074_ (.A1(_03059_),
    .A2(_03148_),
    .B1(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__o31a_1 _08075_ (.A1(_03057_),
    .A2(_03058_),
    .A3(_03148_),
    .B1(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__inv_1 _08076_ (.A(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__nor2_1 _08077_ (.A(_03152_),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__xnor2_1 _08078_ (.A(_03146_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__a21oi_1 _08079_ (.A1(net609),
    .A2(_03158_),
    .B1(_02853_),
    .Y(_03159_));
 sky130_fd_sc_hd__a21o_1 _08080_ (.A1(_00145_),
    .A2(_00138_),
    .B1(_00144_),
    .X(_03160_));
 sky130_fd_sc_hd__a31oi_1 _08081_ (.A1(_00139_),
    .A2(_00145_),
    .A3(_03084_),
    .B1(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__xnor2_1 _08082_ (.A(_00151_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__mux4_2 _08083_ (.A0(\core.CPU_src1_value_a3[18] ),
    .A1(\core.CPU_src1_value_a3[19] ),
    .A2(\core.CPU_src1_value_a3[20] ),
    .A3(\core.CPU_src1_value_a3[21] ),
    .S0(net554),
    .S1(net548),
    .X(_03163_));
 sky130_fd_sc_hd__mux2i_1 _08084_ (.A0(_02983_),
    .A1(_03163_),
    .S(net553),
    .Y(_03164_));
 sky130_fd_sc_hd__mux2i_1 _08085_ (.A0(_02797_),
    .A1(_03164_),
    .S(net478),
    .Y(_03165_));
 sky130_fd_sc_hd__o2bb2ai_1 _08086_ (.A1_N(\core.CPU_is_sll_a3 ),
    .A2_N(_02981_),
    .B1(_02918_),
    .B2(\core.CPU_imm_a3[5] ),
    .Y(_03166_));
 sky130_fd_sc_hd__nand2_1 _08087_ (.A(net478),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__o21ai_0 _08088_ (.A1(_02801_),
    .A2(_03167_),
    .B1(net556),
    .Y(_03168_));
 sky130_fd_sc_hd__a221o_1 _08089_ (.A1(net546),
    .A2(_03162_),
    .B1(_03165_),
    .B2(_02667_),
    .C1(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__nor4_1 _08090_ (.A(_00130_),
    .B(_00136_),
    .C(_00142_),
    .D(_00148_),
    .Y(_03170_));
 sky130_fd_sc_hd__o211ai_1 _08091_ (.A1(_00087_),
    .A2(_02712_),
    .B1(_02782_),
    .C1(_02682_),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _08092_ (.A(_02996_),
    .B(_03170_),
    .Y(_03172_));
 sky130_fd_sc_hd__a21oi_1 _08093_ (.A1(_02806_),
    .A2(_03171_),
    .B1(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__nor2_1 _08094_ (.A(_00142_),
    .B(_00148_),
    .Y(_03174_));
 sky130_fd_sc_hd__a21oi_1 _08095_ (.A1(_03051_),
    .A2(_03174_),
    .B1(_00149_),
    .Y(_03175_));
 sky130_fd_sc_hd__o21ai_0 _08096_ (.A1(_00148_),
    .A2(_03121_),
    .B1(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__a211oi_1 _08097_ (.A1(_02999_),
    .A2(_03170_),
    .B1(_03173_),
    .C1(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__nor2_1 _08098_ (.A(_00053_),
    .B(_02705_),
    .Y(_03178_));
 sky130_fd_sc_hd__or4_1 _08099_ (.A(_00056_),
    .B(_00062_),
    .C(_00070_),
    .D(_00076_),
    .X(_03179_));
 sky130_fd_sc_hd__a21oi_1 _08100_ (.A1(_02704_),
    .A2(_03178_),
    .B1(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__o311a_1 _08101_ (.A1(_02600_),
    .A2(_00062_),
    .A3(_00070_),
    .B1(_02601_),
    .C1(_02602_),
    .X(_03181_));
 sky130_fd_sc_hd__o21bai_1 _08102_ (.A1(_00076_),
    .A2(_03181_),
    .B1_N(_00077_),
    .Y(_03182_));
 sky130_fd_sc_hd__and3_1 _08103_ (.A(_02592_),
    .B(_02610_),
    .C(_02899_),
    .X(_03183_));
 sky130_fd_sc_hd__o2111ai_1 _08104_ (.A1(_03180_),
    .A2(_03182_),
    .B1(_03183_),
    .C1(net438),
    .D1(_03174_),
    .Y(_03184_));
 sky130_fd_sc_hd__nand2_1 _08105_ (.A(net392),
    .B(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__xnor2_1 _08106_ (.A(_00154_),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__a22o_1 _08107_ (.A1(net611),
    .A2(_03162_),
    .B1(_03186_),
    .B2(net476),
    .X(_03187_));
 sky130_fd_sc_hd__a21o_1 _08108_ (.A1(_03159_),
    .A2(_03169_),
    .B1(_03187_),
    .X(_03188_));
 sky130_fd_sc_hd__nor2_1 _08109_ (.A(\core.CPU_dmem_rd_data_a5[21] ),
    .B(net535),
    .Y(_03189_));
 sky130_fd_sc_hd__nor2_1 _08110_ (.A(\core.CPU_reset_a3 ),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__o21ai_1 _08111_ (.A1(net562),
    .A2(_03188_),
    .B1(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__nand3_1 _08113_ (.A(\core.CPU_Xreg_value_a4[10][21] ),
    .B(net550),
    .C(net428),
    .Y(_03193_));
 sky130_fd_sc_hd__o21ai_0 _08114_ (.A1(net428),
    .A2(net356),
    .B1(_03193_),
    .Y(_00765_));
 sky130_fd_sc_hd__nand2_1 _08115_ (.A(\core.CPU_Xreg_value_a4[10][22] ),
    .B(_02563_),
    .Y(_03194_));
 sky130_fd_sc_hd__mux4_2 _08116_ (.A0(\core.CPU_src1_value_a3[19] ),
    .A1(\core.CPU_src1_value_a3[20] ),
    .A2(\core.CPU_src1_value_a3[21] ),
    .A3(\core.CPU_src1_value_a3[22] ),
    .S0(net554),
    .S1(net548),
    .X(_03195_));
 sky130_fd_sc_hd__mux2i_1 _08117_ (.A0(_03010_),
    .A1(_03195_),
    .S(net553),
    .Y(_03196_));
 sky130_fd_sc_hd__nand2_1 _08118_ (.A(_02982_),
    .B(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__o211ai_1 _08119_ (.A1(_02982_),
    .A2(_02838_),
    .B1(_03197_),
    .C1(net478),
    .Y(_03198_));
 sky130_fd_sc_hd__nand3_1 _08120_ (.A(_02982_),
    .B(net480),
    .C(_02835_),
    .Y(_03199_));
 sky130_fd_sc_hd__a21oi_1 _08121_ (.A1(_03198_),
    .A2(_03199_),
    .B1(net475),
    .Y(_03200_));
 sky130_fd_sc_hd__nand2_1 _08122_ (.A(_00145_),
    .B(_00151_),
    .Y(_03201_));
 sky130_fd_sc_hd__a21oi_1 _08123_ (.A1(_00151_),
    .A2(_00144_),
    .B1(_00150_),
    .Y(_03202_));
 sky130_fd_sc_hd__o21ai_0 _08124_ (.A1(_03133_),
    .A2(_03201_),
    .B1(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__a211oi_1 _08125_ (.A1(_02820_),
    .A2(_02822_),
    .B1(_03017_),
    .C1(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__nor2_1 _08126_ (.A(_03130_),
    .B(_03201_),
    .Y(_03205_));
 sky130_fd_sc_hd__o211ai_1 _08127_ (.A1(_02941_),
    .A2(_03015_),
    .B1(_03018_),
    .C1(_03016_),
    .Y(_03206_));
 sky130_fd_sc_hd__a21oi_1 _08128_ (.A1(_03205_),
    .A2(_03206_),
    .B1(_03203_),
    .Y(_03207_));
 sky130_fd_sc_hd__a21oi_1 _08129_ (.A1(_02829_),
    .A2(_03204_),
    .B1(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__xnor2_1 _08130_ (.A(_00157_),
    .B(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__nor2_1 _08131_ (.A(_02540_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__o21bai_1 _08132_ (.A1(_03200_),
    .A2(_03210_),
    .B1_N(_02979_),
    .Y(_03211_));
 sky130_fd_sc_hd__nor3_1 _08133_ (.A(_01127_),
    .B(_01130_),
    .C(_01133_),
    .Y(_03212_));
 sky130_fd_sc_hd__o211ai_1 _08134_ (.A1(_03025_),
    .A2(_03026_),
    .B1(_03111_),
    .C1(_03027_),
    .Y(_03213_));
 sky130_fd_sc_hd__a21o_1 _08135_ (.A1(_00154_),
    .A2(_00147_),
    .B1(_00153_),
    .X(_03214_));
 sky130_fd_sc_hd__a41oi_1 _08136_ (.A1(_00148_),
    .A2(_00154_),
    .A3(_03112_),
    .A4(_03213_),
    .B1(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__a21boi_0 _08137_ (.A1(_02851_),
    .A2(_03212_),
    .B1_N(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__xnor2_1 _08138_ (.A(_00160_),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__nor2_1 _08139_ (.A(net557),
    .B(_03209_),
    .Y(_03218_));
 sky130_fd_sc_hd__a21oi_1 _08140_ (.A1(_00149_),
    .A2(_03146_),
    .B1(_00155_),
    .Y(_03219_));
 sky130_fd_sc_hd__nor2_1 _08141_ (.A(_00148_),
    .B(_00154_),
    .Y(_03220_));
 sky130_fd_sc_hd__o21ai_0 _08142_ (.A1(_00143_),
    .A2(_03120_),
    .B1(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__o2111ai_1 _08143_ (.A1(_03032_),
    .A2(_03033_),
    .B1(_03219_),
    .C1(_03221_),
    .D1(_03037_),
    .Y(_03222_));
 sky130_fd_sc_hd__inv_1 _08144_ (.A(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__nand2_1 _08145_ (.A(_03123_),
    .B(_03220_),
    .Y(_03224_));
 sky130_fd_sc_hd__and3_1 _08146_ (.A(_03219_),
    .B(_03221_),
    .C(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__a21oi_1 _08147_ (.A1(_03035_),
    .A2(_03223_),
    .B1(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__nor3_1 _08148_ (.A(_00160_),
    .B(_02804_),
    .C(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__and3_1 _08149_ (.A(_00160_),
    .B(net476),
    .C(_03226_),
    .X(_03228_));
 sky130_fd_sc_hd__a2111oi_0 _08150_ (.A1(_03127_),
    .A2(_03217_),
    .B1(_03218_),
    .C1(_03227_),
    .D1(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__nor2_1 _08151_ (.A(\core.CPU_dmem_rd_data_a5[22] ),
    .B(net536),
    .Y(_03230_));
 sky130_fd_sc_hd__a31oi_2 _08152_ (.A1(net535),
    .A2(_03211_),
    .A3(net369),
    .B1(net437),
    .Y(_03231_));
 sky130_fd_sc_hd__nand2_1 _08153_ (.A(net429),
    .B(net355),
    .Y(_03232_));
 sky130_fd_sc_hd__a21oi_1 _08154_ (.A1(_03194_),
    .A2(_03232_),
    .B1(net607),
    .Y(_00766_));
 sky130_fd_sc_hd__nand2_1 _08155_ (.A(_00139_),
    .B(_00157_),
    .Y(_03233_));
 sky130_fd_sc_hd__nor2_1 _08156_ (.A(_03201_),
    .B(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__a21o_1 _08157_ (.A1(_00151_),
    .A2(_03160_),
    .B1(_00150_),
    .X(_03235_));
 sky130_fd_sc_hd__a221oi_1 _08158_ (.A1(_03082_),
    .A2(_03234_),
    .B1(_03235_),
    .B2(_00157_),
    .C1(_00156_),
    .Y(_03236_));
 sky130_fd_sc_hd__nand3_1 _08159_ (.A(_02883_),
    .B(_03077_),
    .C(_03234_),
    .Y(_03237_));
 sky130_fd_sc_hd__a21o_1 _08160_ (.A1(net435),
    .A2(_02884_),
    .B1(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__a21boi_0 _08161_ (.A1(_03236_),
    .A2(_03238_),
    .B1_N(_00163_),
    .Y(_03239_));
 sky130_fd_sc_hd__nand3b_1 _08162_ (.A_N(_00163_),
    .B(_03236_),
    .C(_03238_),
    .Y(_03240_));
 sky130_fd_sc_hd__nand3b_1 _08163_ (.A_N(_03239_),
    .B(_03240_),
    .C(net611),
    .Y(_03241_));
 sky130_fd_sc_hd__inv_1 _08164_ (.A(_00148_),
    .Y(_03242_));
 sky130_fd_sc_hd__a21oi_1 _08165_ (.A1(_00143_),
    .A2(_03242_),
    .B1(_00149_),
    .Y(_03243_));
 sky130_fd_sc_hd__inv_1 _08166_ (.A(_00160_),
    .Y(_03244_));
 sky130_fd_sc_hd__nand2_1 _08167_ (.A(_03146_),
    .B(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__a21oi_1 _08168_ (.A1(_00155_),
    .A2(_03244_),
    .B1(_00161_),
    .Y(_03246_));
 sky130_fd_sc_hd__o2111ai_1 _08169_ (.A1(_03243_),
    .A2(_03245_),
    .B1(_03246_),
    .C1(_03050_),
    .D1(_03052_),
    .Y(_03247_));
 sky130_fd_sc_hd__nor2_1 _08170_ (.A(_02901_),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__nor3_1 _08171_ (.A(_00142_),
    .B(_00148_),
    .C(_03245_),
    .Y(_03249_));
 sky130_fd_sc_hd__o21ai_0 _08172_ (.A1(_03243_),
    .A2(_03245_),
    .B1(_03246_),
    .Y(_03250_));
 sky130_fd_sc_hd__o22ai_1 _08173_ (.A1(net438),
    .A2(_03247_),
    .B1(_03249_),
    .B2(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__a21oi_1 _08174_ (.A1(_02904_),
    .A2(_03248_),
    .B1(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__xnor2_1 _08175_ (.A(_00166_),
    .B(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__nand2_1 _08176_ (.A(net480),
    .B(_02892_),
    .Y(_03254_));
 sky130_fd_sc_hd__mux4_2 _08177_ (.A0(\core.CPU_src1_value_a3[20] ),
    .A1(\core.CPU_src1_value_a3[21] ),
    .A2(\core.CPU_src1_value_a3[22] ),
    .A3(\core.CPU_src1_value_a3[23] ),
    .S0(net554),
    .S1(net548),
    .X(_03255_));
 sky130_fd_sc_hd__mux2i_1 _08178_ (.A0(_03068_),
    .A1(_03255_),
    .S(net553),
    .Y(_03256_));
 sky130_fd_sc_hd__nand2_1 _08179_ (.A(net478),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__o21ai_0 _08180_ (.A1(_02894_),
    .A2(_03167_),
    .B1(_02517_),
    .Y(_03258_));
 sky130_fd_sc_hd__a31oi_1 _08181_ (.A1(_02667_),
    .A2(_03254_),
    .A3(_03257_),
    .B1(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__nor2_1 _08182_ (.A(net611),
    .B(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__nor3b_1 _08183_ (.A(_02540_),
    .B(_03239_),
    .C_N(_03240_),
    .Y(_03261_));
 sky130_fd_sc_hd__inv_1 _08184_ (.A(_00147_),
    .Y(_03262_));
 sky130_fd_sc_hd__o21ai_0 _08185_ (.A1(_00142_),
    .A2(_00141_),
    .B1(_00148_),
    .Y(_03263_));
 sky130_fd_sc_hd__nand2_1 _08186_ (.A(_00154_),
    .B(_00160_),
    .Y(_03264_));
 sky130_fd_sc_hd__a21oi_1 _08187_ (.A1(_03262_),
    .A2(_03263_),
    .B1(_03264_),
    .Y(_03265_));
 sky130_fd_sc_hd__o211ai_1 _08188_ (.A1(_02973_),
    .A2(_03057_),
    .B1(_03153_),
    .C1(_03059_),
    .Y(_03266_));
 sky130_fd_sc_hd__a221o_1 _08189_ (.A1(_00160_),
    .A2(_00153_),
    .B1(_03265_),
    .B2(_03266_),
    .C1(_00159_),
    .X(_03267_));
 sky130_fd_sc_hd__nor3_1 _08190_ (.A(_03147_),
    .B(_03148_),
    .C(_03264_),
    .Y(_03268_));
 sky130_fd_sc_hd__nand2_1 _08191_ (.A(_02877_),
    .B(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__a21oi_1 _08192_ (.A1(_02696_),
    .A2(_02874_),
    .B1(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__o21a_1 _08193_ (.A1(_03267_),
    .A2(_03270_),
    .B1(_00166_),
    .X(_03271_));
 sky130_fd_sc_hd__nor3_1 _08194_ (.A(_00166_),
    .B(_03267_),
    .C(_03270_),
    .Y(_03272_));
 sky130_fd_sc_hd__o21ai_0 _08195_ (.A1(_03271_),
    .A2(_03272_),
    .B1(net477),
    .Y(_03273_));
 sky130_fd_sc_hd__o221ai_1 _08196_ (.A1(net555),
    .A2(_03253_),
    .B1(_03260_),
    .B2(_03261_),
    .C1(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__nor2_1 _08197_ (.A(\core.CPU_dmem_rd_data_a5[23] ),
    .B(net536),
    .Y(_03275_));
 sky130_fd_sc_hd__a31oi_2 _08198_ (.A1(net535),
    .A2(_03241_),
    .A3(_03274_),
    .B1(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand2_1 _08199_ (.A(net429),
    .B(net368),
    .Y(_03277_));
 sky130_fd_sc_hd__nand2_1 _08200_ (.A(\core.CPU_Xreg_value_a4[10][23] ),
    .B(net428),
    .Y(_03278_));
 sky130_fd_sc_hd__a21oi_1 _08201_ (.A1(_03277_),
    .A2(_03278_),
    .B1(net606),
    .Y(_00767_));
 sky130_fd_sc_hd__clkinv_1 _08202_ (.A(_00172_),
    .Y(_03279_));
 sky130_fd_sc_hd__a21o_1 _08203_ (.A1(_00166_),
    .A2(_00159_),
    .B1(_00165_),
    .X(_03280_));
 sky130_fd_sc_hd__a31oi_1 _08204_ (.A1(_00160_),
    .A2(_00166_),
    .A3(_03214_),
    .B1(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__inv_1 _08205_ (.A(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__a311oi_1 _08206_ (.A1(net393),
    .A2(_03113_),
    .A3(_03116_),
    .B1(_01136_),
    .C1(_01133_),
    .Y(_03283_));
 sky130_fd_sc_hd__nor4_1 _08207_ (.A(net556),
    .B(_03279_),
    .C(_03282_),
    .D(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__nand3_1 _08208_ (.A(net553),
    .B(net480),
    .C(net479),
    .Y(_03285_));
 sky130_fd_sc_hd__o21ai_0 _08209_ (.A1(net480),
    .A2(_02921_),
    .B1(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hd__mux4_2 _08210_ (.A0(\core.CPU_src1_value_a3[21] ),
    .A1(\core.CPU_src1_value_a3[22] ),
    .A2(\core.CPU_src1_value_a3[23] ),
    .A3(\core.CPU_src1_value_a3[24] ),
    .S0(net554),
    .S1(net548),
    .X(_03287_));
 sky130_fd_sc_hd__mux4_2 _08211_ (.A0(_02743_),
    .A1(_02925_),
    .A2(_03102_),
    .A3(_03287_),
    .S0(net553),
    .S1(net478),
    .X(_03288_));
 sky130_fd_sc_hd__and2_0 _08212_ (.A(_02920_),
    .B(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__a311o_1 _08213_ (.A1(net474),
    .A2(_02929_),
    .A3(_03286_),
    .B1(_03289_),
    .C1(_02853_),
    .X(_03290_));
 sky130_fd_sc_hd__o211ai_1 _08214_ (.A1(_03282_),
    .A2(_03283_),
    .B1(net609),
    .C1(_03279_),
    .Y(_03291_));
 sky130_fd_sc_hd__nor3b_2 _08215_ (.A(_03284_),
    .B(_03290_),
    .C_N(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__nand2_1 _08216_ (.A(_03087_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__o21a_1 _08217_ (.A1(_00157_),
    .A2(_00156_),
    .B1(_00163_),
    .X(_03294_));
 sky130_fd_sc_hd__and2_1 _08218_ (.A(_00145_),
    .B(_00151_),
    .X(_03295_));
 sky130_fd_sc_hd__nand2_1 _08219_ (.A(_03135_),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__o211ai_1 _08220_ (.A1(_02735_),
    .A2(_02737_),
    .B1(_03136_),
    .C1(_03295_),
    .Y(_03297_));
 sky130_fd_sc_hd__nand4b_1 _08221_ (.A_N(_00156_),
    .B(_03202_),
    .C(_03296_),
    .D(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__a21oi_1 _08222_ (.A1(_03294_),
    .A2(_03298_),
    .B1(_00162_),
    .Y(_03299_));
 sky130_fd_sc_hd__xnor2_1 _08223_ (.A(_00169_),
    .B(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__a2bb2o_2 _08224_ (.A1_N(net611),
    .A2_N(_03292_),
    .B1(_03293_),
    .B2(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__inv_1 _08225_ (.A(_00166_),
    .Y(_03302_));
 sky130_fd_sc_hd__nand3_1 _08226_ (.A(_03244_),
    .B(_03302_),
    .C(_03220_),
    .Y(_03303_));
 sky130_fd_sc_hd__o21bai_1 _08227_ (.A1(_00160_),
    .A2(_03219_),
    .B1_N(_00161_),
    .Y(_03304_));
 sky130_fd_sc_hd__a21oi_1 _08228_ (.A1(_03302_),
    .A2(_03304_),
    .B1(_00167_),
    .Y(_03305_));
 sky130_fd_sc_hd__o21ai_0 _08229_ (.A1(_03125_),
    .A2(_03303_),
    .B1(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__xnor2_1 _08230_ (.A(_03279_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__a21oi_1 _08231_ (.A1(net476),
    .A2(_03307_),
    .B1(net562),
    .Y(_03308_));
 sky130_fd_sc_hd__a22oi_4 _08232_ (.A1(\core.CPU_dmem_rd_data_a5[24] ),
    .A2(net562),
    .B1(_03301_),
    .B2(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__o21ai_0 _08234_ (.A1(\core.CPU_Xreg_value_a4[10][24] ),
    .A2(net429),
    .B1(net552),
    .Y(_03311_));
 sky130_fd_sc_hd__a21oi_1 _08235_ (.A1(net429),
    .A2(_03309_),
    .B1(_03311_),
    .Y(_00768_));
 sky130_fd_sc_hd__inv_1 _08237_ (.A(_00178_),
    .Y(_03313_));
 sky130_fd_sc_hd__nand4_1 _08238_ (.A(_00154_),
    .B(_00160_),
    .C(_00166_),
    .D(_00172_),
    .Y(_03314_));
 sky130_fd_sc_hd__o21bai_1 _08239_ (.A1(_03152_),
    .A2(_03156_),
    .B1_N(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__a21oi_1 _08240_ (.A1(_00166_),
    .A2(_00159_),
    .B1(_00165_),
    .Y(_03316_));
 sky130_fd_sc_hd__nand3_1 _08241_ (.A(_00160_),
    .B(_00166_),
    .C(_00153_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21oi_1 _08242_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_03279_),
    .Y(_03318_));
 sky130_fd_sc_hd__nor2_1 _08243_ (.A(_00171_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__nand3_1 _08244_ (.A(_03313_),
    .B(_03315_),
    .C(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__a21o_1 _08245_ (.A1(_03315_),
    .A2(_03319_),
    .B1(_03313_),
    .X(_03321_));
 sky130_fd_sc_hd__nand2_1 _08246_ (.A(net474),
    .B(_02989_),
    .Y(_03322_));
 sky130_fd_sc_hd__nand2_1 _08247_ (.A(net481),
    .B(_03163_),
    .Y(_03323_));
 sky130_fd_sc_hd__mux4_2 _08248_ (.A0(\core.CPU_src1_value_a3[22] ),
    .A1(\core.CPU_src1_value_a3[23] ),
    .A2(\core.CPU_src1_value_a3[24] ),
    .A3(\core.CPU_src1_value_a3[25] ),
    .S0(net554),
    .S1(net548),
    .X(_03324_));
 sky130_fd_sc_hd__nand2_1 _08249_ (.A(net553),
    .B(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__nand3_1 _08250_ (.A(_02982_),
    .B(_03323_),
    .C(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__nand4_1 _08251_ (.A(net478),
    .B(_02929_),
    .C(_03322_),
    .D(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__nand3_1 _08252_ (.A(net480),
    .B(_02929_),
    .C(_02988_),
    .Y(_03328_));
 sky130_fd_sc_hd__nand3_1 _08253_ (.A(net547),
    .B(_03327_),
    .C(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__a31oi_1 _08254_ (.A1(net609),
    .A2(_03320_),
    .A3(_03321_),
    .B1(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__a21o_1 _08255_ (.A1(_00169_),
    .A2(_00162_),
    .B1(_00168_),
    .X(_03331_));
 sky130_fd_sc_hd__nand2_1 _08256_ (.A(_00163_),
    .B(_00169_),
    .Y(_03332_));
 sky130_fd_sc_hd__a21oi_1 _08257_ (.A1(_03236_),
    .A2(_03238_),
    .B1(_03332_),
    .Y(_03333_));
 sky130_fd_sc_hd__nand2b_1 _08259_ (.A_N(_00175_),
    .B(net611),
    .Y(_03335_));
 sky130_fd_sc_hd__o211ai_1 _08260_ (.A1(_03331_),
    .A2(_03333_),
    .B1(net611),
    .C1(_00175_),
    .Y(_03336_));
 sky130_fd_sc_hd__a21o_1 _08261_ (.A1(net392),
    .A2(_03184_),
    .B1(_03245_),
    .X(_03337_));
 sky130_fd_sc_hd__a21oi_1 _08262_ (.A1(_00167_),
    .A2(_03279_),
    .B1(_00173_),
    .Y(_03338_));
 sky130_fd_sc_hd__nand2_1 _08263_ (.A(_03246_),
    .B(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__nor3_1 _08264_ (.A(_03313_),
    .B(_02804_),
    .C(_03339_),
    .Y(_03340_));
 sky130_fd_sc_hd__or2_0 _08265_ (.A(_00166_),
    .B(_00172_),
    .X(_03341_));
 sky130_fd_sc_hd__or3_1 _08266_ (.A(_00178_),
    .B(_02804_),
    .C(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__a211oi_1 _08267_ (.A1(net392),
    .A2(_03184_),
    .B1(_03245_),
    .C1(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__or4_1 _08268_ (.A(_00178_),
    .B(_02804_),
    .C(_03246_),
    .D(_03341_),
    .X(_03344_));
 sky130_fd_sc_hd__nand4_1 _08269_ (.A(_00178_),
    .B(_02864_),
    .C(_03338_),
    .D(_03341_),
    .Y(_03345_));
 sky130_fd_sc_hd__o311ai_0 _08270_ (.A1(_00178_),
    .A2(_02804_),
    .A3(_03338_),
    .B1(_03344_),
    .C1(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__a211oi_1 _08271_ (.A1(_03337_),
    .A2(_03340_),
    .B1(_03343_),
    .C1(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__o311ai_0 _08272_ (.A1(_03331_),
    .A2(_03333_),
    .A3(_03335_),
    .B1(_03336_),
    .C1(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__nor3_1 _08273_ (.A(_00175_),
    .B(_03331_),
    .C(_03333_),
    .Y(_03349_));
 sky130_fd_sc_hd__o21ai_0 _08274_ (.A1(_03331_),
    .A2(_03333_),
    .B1(_00175_),
    .Y(_03350_));
 sky130_fd_sc_hd__nand4b_1 _08275_ (.A_N(_03349_),
    .B(_02915_),
    .C(_03350_),
    .D(_03347_),
    .Y(_03351_));
 sky130_fd_sc_hd__o21ai_0 _08276_ (.A1(_03330_),
    .A2(_03348_),
    .B1(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__mux2i_1 _08277_ (.A0(\core.CPU_dmem_rd_data_a5[25] ),
    .A1(_03352_),
    .S(net535),
    .Y(_03353_));
 sky130_fd_sc_hd__o21ai_0 _08278_ (.A1(\core.CPU_Xreg_value_a4[10][25] ),
    .A2(net429),
    .B1(_02644_),
    .Y(_03354_));
 sky130_fd_sc_hd__a21oi_1 _08279_ (.A1(net429),
    .A2(net354),
    .B1(_03354_),
    .Y(_00769_));
 sky130_fd_sc_hd__nor2_1 _08280_ (.A(\core.CPU_imm_a3[5] ),
    .B(_02918_),
    .Y(_03355_));
 sky130_fd_sc_hd__a21oi_1 _08281_ (.A1(\core.CPU_is_sll_a3 ),
    .A2(_02981_),
    .B1(_03355_),
    .Y(_03356_));
 sky130_fd_sc_hd__mux4_2 _08282_ (.A0(\core.CPU_src1_value_a3[23] ),
    .A1(\core.CPU_src1_value_a3[24] ),
    .A2(\core.CPU_src1_value_a3[25] ),
    .A3(\core.CPU_src1_value_a3[26] ),
    .S0(net554),
    .S1(net548),
    .X(_03357_));
 sky130_fd_sc_hd__mux4_2 _08283_ (.A0(_02833_),
    .A1(_03010_),
    .A2(_03195_),
    .A3(_03357_),
    .S0(net553),
    .S1(net478),
    .X(_03358_));
 sky130_fd_sc_hd__a21oi_1 _08284_ (.A1(_02667_),
    .A2(_03358_),
    .B1(_02979_),
    .Y(_03359_));
 sky130_fd_sc_hd__o21ai_1 _08285_ (.A1(_02589_),
    .A2(_03356_),
    .B1(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__a21o_1 _08286_ (.A1(_00163_),
    .A2(_00156_),
    .B1(_00162_),
    .X(_03361_));
 sky130_fd_sc_hd__a21o_1 _08287_ (.A1(_00169_),
    .A2(_03361_),
    .B1(_00168_),
    .X(_03362_));
 sky130_fd_sc_hd__a21o_1 _08288_ (.A1(_00175_),
    .A2(_03362_),
    .B1(_00174_),
    .X(_03363_));
 sky130_fd_sc_hd__nand4_1 _08289_ (.A(_00157_),
    .B(_00163_),
    .C(_00169_),
    .D(_00175_),
    .Y(_03364_));
 sky130_fd_sc_hd__a211oi_1 _08290_ (.A1(_02829_),
    .A2(_03204_),
    .B1(_03364_),
    .C1(_03207_),
    .Y(_03365_));
 sky130_fd_sc_hd__o21ai_0 _08292_ (.A1(_03363_),
    .A2(_03365_),
    .B1(_00181_),
    .Y(_03367_));
 sky130_fd_sc_hd__or3_1 _08293_ (.A(_00181_),
    .B(_03363_),
    .C(_03365_),
    .X(_03368_));
 sky130_fd_sc_hd__o211ai_1 _08294_ (.A1(net546),
    .A2(_03360_),
    .B1(_03367_),
    .C1(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__nand2_1 _08295_ (.A(net557),
    .B(_03360_),
    .Y(_03370_));
 sky130_fd_sc_hd__a21o_1 _08296_ (.A1(_00172_),
    .A2(_03280_),
    .B1(_00171_),
    .X(_03371_));
 sky130_fd_sc_hd__a21oi_1 _08297_ (.A1(_00178_),
    .A2(_03371_),
    .B1(_00177_),
    .Y(_03372_));
 sky130_fd_sc_hd__o41ai_1 _08298_ (.A1(_03279_),
    .A2(_03313_),
    .A3(_01136_),
    .A4(_03215_),
    .B1(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__a41oi_1 _08299_ (.A1(_00172_),
    .A2(_00178_),
    .A3(_01137_),
    .A4(_02851_),
    .B1(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__nor2b_1 _08300_ (.A(_00166_),
    .B_N(_00161_),
    .Y(_03375_));
 sky130_fd_sc_hd__o21a_1 _08301_ (.A1(_00167_),
    .A2(_03375_),
    .B1(_03279_),
    .X(_03376_));
 sky130_fd_sc_hd__a311oi_1 _08302_ (.A1(_03219_),
    .A2(_03221_),
    .A3(_03224_),
    .B1(_03341_),
    .C1(_00160_),
    .Y(_03377_));
 sky130_fd_sc_hd__o31ai_1 _08303_ (.A1(_00173_),
    .A2(_03376_),
    .A3(_03377_),
    .B1(_03313_),
    .Y(_03378_));
 sky130_fd_sc_hd__nor4_1 _08304_ (.A(_00173_),
    .B(_03034_),
    .C(_03222_),
    .D(_03376_),
    .Y(_03379_));
 sky130_fd_sc_hd__or3_1 _08305_ (.A(_00173_),
    .B(_02857_),
    .C(_03376_),
    .X(_03380_));
 sky130_fd_sc_hd__nor4_1 _08306_ (.A(net427),
    .B(_02861_),
    .C(_03222_),
    .D(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__inv_1 _08307_ (.A(_00179_),
    .Y(_03382_));
 sky130_fd_sc_hd__o31ai_1 _08308_ (.A1(_03378_),
    .A2(_03379_),
    .A3(_03381_),
    .B1(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__o221ai_1 _08310_ (.A1(_02994_),
    .A2(_03374_),
    .B1(_03383_),
    .B2(_02804_),
    .C1(_00184_),
    .Y(_03385_));
 sky130_fd_sc_hd__a221o_1 _08311_ (.A1(_03127_),
    .A2(_03374_),
    .B1(_03383_),
    .B2(net476),
    .C1(_00184_),
    .X(_03386_));
 sky130_fd_sc_hd__a22o_1 _08312_ (.A1(_03369_),
    .A2(_03370_),
    .B1(_03385_),
    .B2(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__nor2_1 _08313_ (.A(_01114_),
    .B(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__a21oi_2 _08314_ (.A1(\core.CPU_dmem_rd_data_a5[26] ),
    .A2(_01114_),
    .B1(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__o21ai_0 _08315_ (.A1(\core.CPU_Xreg_value_a4[10][26] ),
    .A2(net429),
    .B1(net551),
    .Y(_03390_));
 sky130_fd_sc_hd__a21oi_1 _08316_ (.A1(net429),
    .A2(_03389_),
    .B1(_03390_),
    .Y(_00770_));
 sky130_fd_sc_hd__inv_1 _08317_ (.A(_00029_),
    .Y(_03391_));
 sky130_fd_sc_hd__a21oi_1 _08318_ (.A1(_00172_),
    .A2(_00165_),
    .B1(_00171_),
    .Y(_03392_));
 sky130_fd_sc_hd__o21bai_1 _08319_ (.A1(_03313_),
    .A2(_03392_),
    .B1_N(_00177_),
    .Y(_03393_));
 sky130_fd_sc_hd__a21oi_1 _08320_ (.A1(_00184_),
    .A2(_03393_),
    .B1(_00183_),
    .Y(_03394_));
 sky130_fd_sc_hd__nand3_1 _08321_ (.A(_00166_),
    .B(_01157_),
    .C(_03267_),
    .Y(_03395_));
 sky130_fd_sc_hd__nand3_1 _08322_ (.A(_00166_),
    .B(_01157_),
    .C(_03270_),
    .Y(_03396_));
 sky130_fd_sc_hd__a31oi_1 _08323_ (.A1(_03394_),
    .A2(_03395_),
    .A3(_03396_),
    .B1(_02609_),
    .Y(_03397_));
 sky130_fd_sc_hd__nor3_1 _08324_ (.A(_00178_),
    .B(_00184_),
    .C(_03341_),
    .Y(_03398_));
 sky130_fd_sc_hd__nand2_1 _08325_ (.A(_03252_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__inv_1 _08326_ (.A(_00184_),
    .Y(_03400_));
 sky130_fd_sc_hd__o21ai_0 _08327_ (.A1(_00178_),
    .A2(_03338_),
    .B1(_03382_),
    .Y(_03401_));
 sky130_fd_sc_hd__a21oi_1 _08328_ (.A1(_03400_),
    .A2(_03401_),
    .B1(_00185_),
    .Y(_03402_));
 sky130_fd_sc_hd__and3_1 _08329_ (.A(net612),
    .B(_03399_),
    .C(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__a21oi_1 _08330_ (.A1(_03399_),
    .A2(_03402_),
    .B1(net555),
    .Y(_03404_));
 sky130_fd_sc_hd__o211ai_1 _08331_ (.A1(_03267_),
    .A2(_03270_),
    .B1(_00166_),
    .C1(_01157_),
    .Y(_03405_));
 sky130_fd_sc_hd__a31o_2 _08332_ (.A1(net477),
    .A2(_03394_),
    .A3(_03405_),
    .B1(_00029_),
    .X(_03406_));
 sky130_fd_sc_hd__o32ai_1 _08333_ (.A1(_03391_),
    .A2(_03397_),
    .A3(_03403_),
    .B1(_03404_),
    .B2(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand4_1 _08334_ (.A(_00163_),
    .B(_00169_),
    .C(_00175_),
    .D(_00181_),
    .Y(_03408_));
 sky130_fd_sc_hd__nand3_1 _08335_ (.A(_00175_),
    .B(_00181_),
    .C(_03331_),
    .Y(_03409_));
 sky130_fd_sc_hd__a21oi_1 _08336_ (.A1(_00181_),
    .A2(_00174_),
    .B1(_00180_),
    .Y(_03410_));
 sky130_fd_sc_hd__nand2_1 _08337_ (.A(_03409_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__o21bai_1 _08338_ (.A1(_03236_),
    .A2(_03408_),
    .B1_N(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__nor3_1 _08339_ (.A(_03076_),
    .B(_03201_),
    .C(_03233_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand2_1 _08340_ (.A(_00175_),
    .B(_00181_),
    .Y(_03414_));
 sky130_fd_sc_hd__nor3_1 _08341_ (.A(_02966_),
    .B(_03332_),
    .C(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand3_1 _08342_ (.A(_02883_),
    .B(_03413_),
    .C(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__a21oi_1 _08343_ (.A1(net435),
    .A2(_02884_),
    .B1(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__or3_1 _08344_ (.A(_00187_),
    .B(_03412_),
    .C(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__o21ai_0 _08345_ (.A1(_03412_),
    .A2(_03417_),
    .B1(_00187_),
    .Y(_03419_));
 sky130_fd_sc_hd__o2111ai_1 _08346_ (.A1(net611),
    .A2(net367),
    .B1(_03418_),
    .C1(_03419_),
    .D1(_02794_),
    .Y(_03420_));
 sky130_fd_sc_hd__a31oi_1 _08348_ (.A1(_02674_),
    .A2(_02678_),
    .A3(_03166_),
    .B1(_02539_),
    .Y(_03422_));
 sky130_fd_sc_hd__nor2_1 _08349_ (.A(net611),
    .B(_02525_),
    .Y(_03423_));
 sky130_fd_sc_hd__mux2i_1 _08350_ (.A0(\core.CPU_src1_value_a3[25] ),
    .A1(\core.CPU_src1_value_a3[27] ),
    .S(net548),
    .Y(_03424_));
 sky130_fd_sc_hd__and2_1 _08351_ (.A(\core.CPU_src1_value_a3[24] ),
    .B(_02577_),
    .X(_03425_));
 sky130_fd_sc_hd__a211oi_1 _08352_ (.A1(\core.CPU_src1_value_a3[26] ),
    .A2(net548),
    .B1(_03425_),
    .C1(net554),
    .Y(_03426_));
 sky130_fd_sc_hd__a21oi_1 _08353_ (.A1(net554),
    .A2(_03424_),
    .B1(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__mux4_2 _08354_ (.A0(_02891_),
    .A1(_03068_),
    .A2(_03255_),
    .A3(_03427_),
    .S0(net553),
    .S1(net478),
    .X(_03428_));
 sky130_fd_sc_hd__nand2_1 _08355_ (.A(_03423_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__o21ai_0 _08356_ (.A1(net611),
    .A2(_03422_),
    .B1(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__nand2_1 _08357_ (.A(net367),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__nor2_1 _08360_ (.A(_01114_),
    .B(net428),
    .Y(_03434_));
 sky130_fd_sc_hd__nor2_1 _08361_ (.A(\core.CPU_dmem_rd_data_a5[27] ),
    .B(net536),
    .Y(_03435_));
 sky130_fd_sc_hd__nand2_1 _08362_ (.A(net429),
    .B(net436),
    .Y(_03436_));
 sky130_fd_sc_hd__o21ai_0 _08363_ (.A1(\core.CPU_Xreg_value_a4[10][27] ),
    .A2(net429),
    .B1(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__a311oi_1 _08365_ (.A1(net353),
    .A2(_03431_),
    .A3(_03434_),
    .B1(_03437_),
    .C1(net606),
    .Y(_00771_));
 sky130_fd_sc_hd__inv_1 _08366_ (.A(_00025_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand4_1 _08367_ (.A(_03391_),
    .B(_03279_),
    .C(_03313_),
    .D(_03400_),
    .Y(_03440_));
 sky130_fd_sc_hd__a21oi_1 _08368_ (.A1(_00173_),
    .A2(_03313_),
    .B1(_00179_),
    .Y(_03441_));
 sky130_fd_sc_hd__nor2_1 _08369_ (.A(_00184_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__o21ai_0 _08370_ (.A1(_00185_),
    .A2(_03442_),
    .B1(_03391_),
    .Y(_03443_));
 sky130_fd_sc_hd__inv_1 _08371_ (.A(_00030_),
    .Y(_03444_));
 sky130_fd_sc_hd__o211ai_1 _08372_ (.A1(_03305_),
    .A2(_03440_),
    .B1(_03443_),
    .C1(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__a211oi_1 _08373_ (.A1(_03122_),
    .A2(_03124_),
    .B1(_03303_),
    .C1(_03440_),
    .Y(_03446_));
 sky130_fd_sc_hd__nor4_1 _08374_ (.A(_03439_),
    .B(net555),
    .C(_03445_),
    .D(_03446_),
    .Y(_03447_));
 sky130_fd_sc_hd__nor2_1 _08375_ (.A(_03439_),
    .B(_02609_),
    .Y(_03448_));
 sky130_fd_sc_hd__nor2_1 _08376_ (.A(_00025_),
    .B(_02609_),
    .Y(_03449_));
 sky130_fd_sc_hd__a21oi_1 _08377_ (.A1(_00178_),
    .A2(_00171_),
    .B1(_00177_),
    .Y(_03450_));
 sky130_fd_sc_hd__o21bai_1 _08378_ (.A1(_03400_),
    .A2(_03450_),
    .B1_N(_00183_),
    .Y(_03451_));
 sky130_fd_sc_hd__a21oi_1 _08379_ (.A1(_00029_),
    .A2(_03451_),
    .B1(_00028_),
    .Y(_03452_));
 sky130_fd_sc_hd__o21ai_0 _08380_ (.A1(_01159_),
    .A2(_03281_),
    .B1(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__a31oi_1 _08381_ (.A1(_00029_),
    .A2(_01157_),
    .A3(_03283_),
    .B1(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__mux2i_1 _08382_ (.A0(_03448_),
    .A1(_03449_),
    .S(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__o211ai_1 _08383_ (.A1(_03445_),
    .A2(_03446_),
    .B1(_03439_),
    .C1(net612),
    .Y(_03456_));
 sky130_fd_sc_hd__nand3b_1 _08384_ (.A_N(_03447_),
    .B(_03455_),
    .C(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__nor2_1 _08385_ (.A(_00187_),
    .B(_00186_),
    .Y(_03458_));
 sky130_fd_sc_hd__nor3_1 _08386_ (.A(_00181_),
    .B(_00180_),
    .C(_00186_),
    .Y(_03459_));
 sky130_fd_sc_hd__nor2_1 _08387_ (.A(_03458_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__o41ai_1 _08388_ (.A1(_00180_),
    .A2(_00186_),
    .A3(_03363_),
    .A4(_03365_),
    .B1(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__xnor2_1 _08389_ (.A(_00189_),
    .B(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__nand2_1 _08390_ (.A(net480),
    .B(_03103_),
    .Y(_03463_));
 sky130_fd_sc_hd__nand2_1 _08391_ (.A(net481),
    .B(_03287_),
    .Y(_03464_));
 sky130_fd_sc_hd__mux2i_1 _08392_ (.A0(\core.CPU_src1_value_a3[26] ),
    .A1(\core.CPU_src1_value_a3[28] ),
    .S(net548),
    .Y(_03465_));
 sky130_fd_sc_hd__mux2i_1 _08393_ (.A0(_03424_),
    .A1(_03465_),
    .S(net554),
    .Y(_03466_));
 sky130_fd_sc_hd__nand2_1 _08394_ (.A(net553),
    .B(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__nand3_1 _08395_ (.A(net478),
    .B(_03464_),
    .C(_03467_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand2_1 _08396_ (.A(net557),
    .B(_02539_),
    .Y(_03469_));
 sky130_fd_sc_hd__o31ai_1 _08397_ (.A1(net611),
    .A2(_02750_),
    .A3(_03356_),
    .B1(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__a31oi_1 _08398_ (.A1(_03423_),
    .A2(_03463_),
    .A3(_03468_),
    .B1(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__a21boi_0 _08399_ (.A1(net546),
    .A2(_03462_),
    .B1_N(net391),
    .Y(_03472_));
 sky130_fd_sc_hd__a21oi_1 _08400_ (.A1(net611),
    .A2(_03462_),
    .B1(_01114_),
    .Y(_03473_));
 sky130_fd_sc_hd__o21ai_1 _08401_ (.A1(_03457_),
    .A2(_03472_),
    .B1(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__nand2b_1 _08402_ (.A_N(\core.CPU_dmem_rd_data_a5[28] ),
    .B(_01114_),
    .Y(_03475_));
 sky130_fd_sc_hd__nand3_1 _08403_ (.A(net429),
    .B(_03474_),
    .C(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_1 _08404_ (.A(\core.CPU_Xreg_value_a4[10][28] ),
    .B(net428),
    .Y(_03477_));
 sky130_fd_sc_hd__a21oi_1 _08405_ (.A1(_03476_),
    .A2(_03477_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_00772_));
 sky130_fd_sc_hd__a21boi_0 _08406_ (.A1(_03316_),
    .A2(_03317_),
    .B1_N(_01157_),
    .Y(_03478_));
 sky130_fd_sc_hd__nor3_1 _08407_ (.A(_00029_),
    .B(_00024_),
    .C(_00028_),
    .Y(_03479_));
 sky130_fd_sc_hd__nor2_1 _08408_ (.A(_00025_),
    .B(_00024_),
    .Y(_03480_));
 sky130_fd_sc_hd__nor2_1 _08409_ (.A(_03479_),
    .B(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__o41ai_1 _08410_ (.A1(_00024_),
    .A2(_00028_),
    .A3(_03451_),
    .A4(_03478_),
    .B1(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__nand2_1 _08411_ (.A(_03155_),
    .B(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__nand4_1 _08412_ (.A(_00025_),
    .B(_00029_),
    .C(_00178_),
    .D(_00184_),
    .Y(_03484_));
 sky130_fd_sc_hd__o21ai_0 _08413_ (.A1(_03314_),
    .A2(_03484_),
    .B1(_03482_),
    .Y(_03485_));
 sky130_fd_sc_hd__o21ai_0 _08414_ (.A1(_03152_),
    .A2(_03483_),
    .B1(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__nor2_1 _08415_ (.A(_00194_),
    .B(_02609_),
    .Y(_03487_));
 sky130_fd_sc_hd__o2111a_1 _08416_ (.A1(_03152_),
    .A2(_03483_),
    .B1(_03485_),
    .C1(_00194_),
    .D1(net477),
    .X(_03488_));
 sky130_fd_sc_hd__a21oi_1 _08417_ (.A1(_03486_),
    .A2(_03487_),
    .B1(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__nor2_1 _08418_ (.A(_00179_),
    .B(_00185_),
    .Y(_03490_));
 sky130_fd_sc_hd__o211ai_1 _08419_ (.A1(_03246_),
    .A2(_03341_),
    .B1(_03490_),
    .C1(_03338_),
    .Y(_03491_));
 sky130_fd_sc_hd__a21oi_1 _08420_ (.A1(_00178_),
    .A2(_03382_),
    .B1(_00184_),
    .Y(_03492_));
 sky130_fd_sc_hd__nor2_1 _08421_ (.A(_00025_),
    .B(_00029_),
    .Y(_03493_));
 sky130_fd_sc_hd__o21a_1 _08422_ (.A1(_00185_),
    .A2(_03492_),
    .B1(_03493_),
    .X(_03494_));
 sky130_fd_sc_hd__a221o_1 _08423_ (.A1(_03439_),
    .A2(_00030_),
    .B1(_03491_),
    .B2(_03494_),
    .C1(_00026_),
    .X(_03495_));
 sky130_fd_sc_hd__nand2_1 _08424_ (.A(net612),
    .B(_00194_),
    .Y(_03496_));
 sky130_fd_sc_hd__nor2_1 _08425_ (.A(_03495_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__nand2_1 _08426_ (.A(_03398_),
    .B(_03493_),
    .Y(_03498_));
 sky130_fd_sc_hd__nand3_1 _08427_ (.A(net612),
    .B(_00194_),
    .C(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__nand2b_1 _08428_ (.A_N(_00194_),
    .B(net612),
    .Y(_03500_));
 sky130_fd_sc_hd__mux2i_1 _08429_ (.A0(_03499_),
    .A1(_03500_),
    .S(_03495_),
    .Y(_03501_));
 sky130_fd_sc_hd__a31oi_1 _08430_ (.A1(net392),
    .A2(_03184_),
    .A3(_03497_),
    .B1(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__nor3_1 _08431_ (.A(_03245_),
    .B(_03498_),
    .C(_03500_),
    .Y(_03503_));
 sky130_fd_sc_hd__nor3b_1 _08432_ (.A(_03495_),
    .B(_03496_),
    .C_N(_03245_),
    .Y(_03504_));
 sky130_fd_sc_hd__a21oi_1 _08433_ (.A1(_03185_),
    .A2(_03503_),
    .B1(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__a31oi_1 _08434_ (.A1(_03489_),
    .A2(_03502_),
    .A3(_03505_),
    .B1(net611),
    .Y(_03506_));
 sky130_fd_sc_hd__nand2_1 _08435_ (.A(_00187_),
    .B(_00189_),
    .Y(_03507_));
 sky130_fd_sc_hd__a211oi_1 _08436_ (.A1(_03236_),
    .A2(_03238_),
    .B1(_03408_),
    .C1(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__a21oi_1 _08437_ (.A1(_00187_),
    .A2(_03411_),
    .B1(_00186_),
    .Y(_03509_));
 sky130_fd_sc_hd__nor2b_1 _08438_ (.A(_03509_),
    .B_N(_00189_),
    .Y(_03510_));
 sky130_fd_sc_hd__or4_1 _08439_ (.A(_00191_),
    .B(_00188_),
    .C(_03508_),
    .D(_03510_),
    .X(_03511_));
 sky130_fd_sc_hd__o31ai_1 _08440_ (.A1(_00188_),
    .A2(_03508_),
    .A3(_03510_),
    .B1(_00191_),
    .Y(_03512_));
 sky130_fd_sc_hd__nand2_1 _08441_ (.A(net480),
    .B(_03164_),
    .Y(_03513_));
 sky130_fd_sc_hd__nand2_1 _08442_ (.A(net481),
    .B(_03324_),
    .Y(_03514_));
 sky130_fd_sc_hd__mux4_2 _08443_ (.A0(\core.CPU_src1_value_a3[26] ),
    .A1(\core.CPU_src1_value_a3[27] ),
    .A2(\core.CPU_src1_value_a3[28] ),
    .A3(\core.CPU_src1_value_a3[29] ),
    .S0(net554),
    .S1(net548),
    .X(_03515_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(net553),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand3_1 _08445_ (.A(net478),
    .B(_03514_),
    .C(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__a31oi_1 _08446_ (.A1(_02667_),
    .A2(_03513_),
    .A3(_03517_),
    .B1(_02539_),
    .Y(_03518_));
 sky130_fd_sc_hd__o21ai_0 _08447_ (.A1(_02802_),
    .A2(_03356_),
    .B1(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__a32oi_1 _08448_ (.A1(_02794_),
    .A2(_03511_),
    .A3(_03512_),
    .B1(_03519_),
    .B2(net557),
    .Y(_03520_));
 sky130_fd_sc_hd__nand2_1 _08449_ (.A(\core.CPU_dmem_rd_data_a5[29] ),
    .B(net562),
    .Y(_03521_));
 sky130_fd_sc_hd__o31ai_1 _08450_ (.A1(_01114_),
    .A2(_03506_),
    .A3(_03520_),
    .B1(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__nand2_1 _08451_ (.A(net549),
    .B(net366),
    .Y(_03523_));
 sky130_fd_sc_hd__nand3_1 _08453_ (.A(\core.CPU_Xreg_value_a4[10][29] ),
    .B(net549),
    .C(net428),
    .Y(_03525_));
 sky130_fd_sc_hd__o21ai_0 _08454_ (.A1(net428),
    .A2(_03523_),
    .B1(_03525_),
    .Y(_00773_));
 sky130_fd_sc_hd__xor2_1 _08455_ (.A(_00008_),
    .B(_00040_),
    .X(_03526_));
 sky130_fd_sc_hd__xnor2_1 _08456_ (.A(_00001_),
    .B(\core.CPU_src1_value_a3[2] ),
    .Y(_03527_));
 sky130_fd_sc_hd__nor2_1 _08457_ (.A(_02540_),
    .B(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__a211o_1 _08458_ (.A1(_02530_),
    .A2(_02586_),
    .B1(_03528_),
    .C1(net609),
    .X(_03529_));
 sky130_fd_sc_hd__nor2b_1 _08459_ (.A(_00040_),
    .B_N(_00005_),
    .Y(_03530_));
 sky130_fd_sc_hd__o21ai_0 _08460_ (.A1(_02611_),
    .A2(_03530_),
    .B1(net609),
    .Y(_03531_));
 sky130_fd_sc_hd__a21oi_1 _08461_ (.A1(_03529_),
    .A2(_03531_),
    .B1(net612),
    .Y(_03532_));
 sky130_fd_sc_hd__a21oi_1 _08462_ (.A1(net612),
    .A2(_03526_),
    .B1(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_1 _08463_ (.A(net611),
    .B(_03527_),
    .Y(_03534_));
 sky130_fd_sc_hd__o21ai_0 _08464_ (.A1(net611),
    .A2(_03533_),
    .B1(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__nand2_1 _08465_ (.A(\core.CPU_dmem_rd_data_a5[2] ),
    .B(net562),
    .Y(_03536_));
 sky130_fd_sc_hd__o21ai_2 _08466_ (.A1(net562),
    .A2(_03535_),
    .B1(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__nor2_1 _08468_ (.A(_02563_),
    .B(net373),
    .Y(_03539_));
 sky130_fd_sc_hd__o21ai_0 _08470_ (.A1(\core.CPU_Xreg_value_a4[10][2] ),
    .A2(_02558_),
    .B1(_02644_),
    .Y(_03541_));
 sky130_fd_sc_hd__nor2_1 _08471_ (.A(_03539_),
    .B(_03541_),
    .Y(_00774_));
 sky130_fd_sc_hd__nor2_1 _08472_ (.A(_00184_),
    .B(_00194_),
    .Y(_03542_));
 sky130_fd_sc_hd__a21oi_1 _08473_ (.A1(_03391_),
    .A2(_00185_),
    .B1(_00030_),
    .Y(_03543_));
 sky130_fd_sc_hd__nor2_1 _08474_ (.A(_00025_),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__nor2_1 _08475_ (.A(_00026_),
    .B(_03544_),
    .Y(_03545_));
 sky130_fd_sc_hd__nor2_1 _08476_ (.A(_00194_),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__a311oi_1 _08477_ (.A1(_03383_),
    .A2(_03493_),
    .A3(_03542_),
    .B1(_03546_),
    .C1(_00195_),
    .Y(_03547_));
 sky130_fd_sc_hd__xnor2_1 _08478_ (.A(_00200_),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__nand4_1 _08479_ (.A(_00025_),
    .B(_00029_),
    .C(_00184_),
    .D(_00194_),
    .Y(_03549_));
 sky130_fd_sc_hd__a21oi_1 _08480_ (.A1(_00029_),
    .A2(_00183_),
    .B1(_00028_),
    .Y(_03550_));
 sky130_fd_sc_hd__nor2b_1 _08481_ (.A(_03550_),
    .B_N(_00025_),
    .Y(_03551_));
 sky130_fd_sc_hd__o21ai_0 _08482_ (.A1(_00024_),
    .A2(_03551_),
    .B1(_00194_),
    .Y(_03552_));
 sky130_fd_sc_hd__nand2b_1 _08483_ (.A_N(_00193_),
    .B(_03552_),
    .Y(_03553_));
 sky130_fd_sc_hd__nor2_1 _08484_ (.A(_00200_),
    .B(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__nand2_1 _08485_ (.A(_03549_),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__nand2_1 _08486_ (.A(_00200_),
    .B(_03553_),
    .Y(_03556_));
 sky130_fd_sc_hd__nor3_1 _08487_ (.A(_03391_),
    .B(_03400_),
    .C(_01163_),
    .Y(_03557_));
 sky130_fd_sc_hd__mux2i_1 _08488_ (.A0(_03557_),
    .A1(_03554_),
    .S(_03374_),
    .Y(_03558_));
 sky130_fd_sc_hd__a31oi_1 _08489_ (.A1(_03555_),
    .A2(_03556_),
    .A3(_03558_),
    .B1(_02609_),
    .Y(_03559_));
 sky130_fd_sc_hd__and3_1 _08490_ (.A(_00187_),
    .B(_00189_),
    .C(_00191_),
    .X(_03560_));
 sky130_fd_sc_hd__a2111o_1 _08491_ (.A1(_00181_),
    .A2(_00174_),
    .B1(_00180_),
    .C1(_00186_),
    .D1(_00190_),
    .X(_03561_));
 sky130_fd_sc_hd__a31oi_1 _08492_ (.A1(_00175_),
    .A2(_00181_),
    .A3(_03362_),
    .B1(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__nand2_1 _08493_ (.A(_00189_),
    .B(_00191_),
    .Y(_03563_));
 sky130_fd_sc_hd__a21oi_1 _08494_ (.A1(_00191_),
    .A2(_00188_),
    .B1(_00190_),
    .Y(_03564_));
 sky130_fd_sc_hd__o31ai_1 _08495_ (.A1(_03458_),
    .A2(_03562_),
    .A3(_03563_),
    .B1(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__a31oi_1 _08496_ (.A1(_00181_),
    .A2(_03365_),
    .A3(_03560_),
    .B1(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__xnor2_1 _08497_ (.A(_00197_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__nor2_1 _08498_ (.A(net611),
    .B(_02540_),
    .Y(_03568_));
 sky130_fd_sc_hd__nand2_1 _08499_ (.A(net481),
    .B(_03357_),
    .Y(_03569_));
 sky130_fd_sc_hd__mux4_2 _08500_ (.A0(\core.CPU_src1_value_a3[27] ),
    .A1(\core.CPU_src1_value_a3[28] ),
    .A2(\core.CPU_src1_value_a3[29] ),
    .A3(\core.CPU_src1_value_a3[30] ),
    .S0(net554),
    .S1(net548),
    .X(_03570_));
 sky130_fd_sc_hd__nand2_1 _08501_ (.A(net553),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__and3_1 _08502_ (.A(net478),
    .B(_03569_),
    .C(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__a211oi_1 _08503_ (.A1(net480),
    .A2(_03196_),
    .B1(_03572_),
    .C1(_02525_),
    .Y(_03573_));
 sky130_fd_sc_hd__a211o_1 _08504_ (.A1(_02839_),
    .A2(_03166_),
    .B1(_03573_),
    .C1(_02539_),
    .X(_03574_));
 sky130_fd_sc_hd__a22oi_1 _08505_ (.A1(_03567_),
    .A2(_03568_),
    .B1(_03574_),
    .B2(net557),
    .Y(_03575_));
 sky130_fd_sc_hd__a211oi_1 _08506_ (.A1(net612),
    .A2(_03548_),
    .B1(_03559_),
    .C1(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__nand3_1 _08507_ (.A(net611),
    .B(net535),
    .C(_03567_),
    .Y(_03577_));
 sky130_fd_sc_hd__nand2_1 _08508_ (.A(\core.CPU_dmem_rd_data_a5[30] ),
    .B(net562),
    .Y(_03578_));
 sky130_fd_sc_hd__nand2_1 _08509_ (.A(_03577_),
    .B(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__a21oi_1 _08510_ (.A1(net535),
    .A2(_03576_),
    .B1(_03579_),
    .Y(_03580_));
 sky130_fd_sc_hd__o21ai_0 _08511_ (.A1(\core.CPU_Xreg_value_a4[10][30] ),
    .A2(net429),
    .B1(_02644_),
    .Y(_03581_));
 sky130_fd_sc_hd__a21oi_1 _08512_ (.A1(net429),
    .A2(net345),
    .B1(_03581_),
    .Y(_00775_));
 sky130_fd_sc_hd__nand4_1 _08513_ (.A(_00025_),
    .B(_00029_),
    .C(_00194_),
    .D(_00200_),
    .Y(_03582_));
 sky130_fd_sc_hd__nor3_1 _08514_ (.A(net556),
    .B(_01155_),
    .C(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__xnor2_1 _08515_ (.A(net585),
    .B(\core.CPU_src1_value_a3[31] ),
    .Y(_03584_));
 sky130_fd_sc_hd__a21o_1 _08516_ (.A1(_00025_),
    .A2(_00028_),
    .B1(_00024_),
    .X(_03585_));
 sky130_fd_sc_hd__a21o_1 _08517_ (.A1(_00194_),
    .A2(_03585_),
    .B1(_00193_),
    .X(_03586_));
 sky130_fd_sc_hd__a21oi_1 _08518_ (.A1(_00200_),
    .A2(_03586_),
    .B1(_00199_),
    .Y(_03587_));
 sky130_fd_sc_hd__nand2_1 _08519_ (.A(_03394_),
    .B(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__nor3_1 _08520_ (.A(net556),
    .B(_03584_),
    .C(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__mux2i_1 _08521_ (.A0(_03583_),
    .A1(_03589_),
    .S(_03405_),
    .Y(_03590_));
 sky130_fd_sc_hd__mux4_2 _08522_ (.A0(\core.CPU_src1_value_a3[28] ),
    .A1(\core.CPU_src1_value_a3[29] ),
    .A2(\core.CPU_src1_value_a3[30] ),
    .A3(\core.CPU_src1_value_a3[31] ),
    .S0(net554),
    .S1(net548),
    .X(_03591_));
 sky130_fd_sc_hd__nor3_1 _08523_ (.A(net553),
    .B(_02525_),
    .C(net480),
    .Y(_03592_));
 sky130_fd_sc_hd__a22oi_1 _08524_ (.A1(net441),
    .A2(_03591_),
    .B1(_03592_),
    .B2(_03427_),
    .Y(_03593_));
 sky130_fd_sc_hd__o22ai_1 _08525_ (.A1(_02894_),
    .A2(_03356_),
    .B1(_03256_),
    .B2(_02525_),
    .Y(_03594_));
 sky130_fd_sc_hd__nand2_1 _08526_ (.A(net480),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__o2111ai_1 _08527_ (.A1(_02892_),
    .A2(_03167_),
    .B1(_03593_),
    .C1(_03595_),
    .D1(net556),
    .Y(_03596_));
 sky130_fd_sc_hd__o21a_1 _08528_ (.A1(_03394_),
    .A2(_03582_),
    .B1(_03587_),
    .X(_03597_));
 sky130_fd_sc_hd__nand3_1 _08529_ (.A(_01155_),
    .B(_03587_),
    .C(_03582_),
    .Y(_03598_));
 sky130_fd_sc_hd__o21ai_0 _08530_ (.A1(_01155_),
    .A2(_03597_),
    .B1(_03598_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand2_1 _08531_ (.A(net609),
    .B(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__a31o_2 _08532_ (.A1(_03590_),
    .A2(_03596_),
    .A3(_03600_),
    .B1(_02853_),
    .X(_03601_));
 sky130_fd_sc_hd__xnor2_1 _08533_ (.A(\core.CPU_src1_value_a3[31] ),
    .B(net613),
    .Y(_03602_));
 sky130_fd_sc_hd__a21o_1 _08534_ (.A1(_00189_),
    .A2(_00186_),
    .B1(_00188_),
    .X(_03603_));
 sky130_fd_sc_hd__a211o_1 _08535_ (.A1(_00191_),
    .A2(_03603_),
    .B1(_00196_),
    .C1(_00190_),
    .X(_03604_));
 sky130_fd_sc_hd__o22a_1 _08536_ (.A1(_00197_),
    .A2(_00196_),
    .B1(_03560_),
    .B2(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__o31ai_1 _08537_ (.A1(_03412_),
    .A2(_03417_),
    .A3(_03604_),
    .B1(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__xnor2_1 _08538_ (.A(_03602_),
    .B(_03606_),
    .Y(_03607_));
 sky130_fd_sc_hd__nand2_1 _08539_ (.A(net611),
    .B(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__o21ai_0 _08540_ (.A1(_03087_),
    .A2(_03607_),
    .B1(net535),
    .Y(_03609_));
 sky130_fd_sc_hd__a21oi_1 _08541_ (.A1(_03601_),
    .A2(_03608_),
    .B1(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__nor2_1 _08543_ (.A(_00201_),
    .B(_01155_),
    .Y(_03612_));
 sky130_fd_sc_hd__nor2_1 _08544_ (.A(_00200_),
    .B(_03584_),
    .Y(_03613_));
 sky130_fd_sc_hd__nor2_1 _08545_ (.A(_00194_),
    .B(_03498_),
    .Y(_03614_));
 sky130_fd_sc_hd__inv_1 _08546_ (.A(_00026_),
    .Y(_03615_));
 sky130_fd_sc_hd__o211ai_1 _08547_ (.A1(_00029_),
    .A2(_03402_),
    .B1(_03615_),
    .C1(_03444_),
    .Y(_03616_));
 sky130_fd_sc_hd__a21oi_1 _08548_ (.A1(_00025_),
    .A2(_03615_),
    .B1(_00194_),
    .Y(_03617_));
 sky130_fd_sc_hd__a221o_1 _08549_ (.A1(_03252_),
    .A2(_03614_),
    .B1(_03616_),
    .B2(_03617_),
    .C1(_00195_),
    .X(_03618_));
 sky130_fd_sc_hd__mux2i_1 _08550_ (.A0(_03612_),
    .A1(_03613_),
    .S(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__nand2_1 _08551_ (.A(_00201_),
    .B(_01155_),
    .Y(_03620_));
 sky130_fd_sc_hd__nand2_1 _08552_ (.A(net535),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__a21oi_1 _08553_ (.A1(_00200_),
    .A2(_03612_),
    .B1(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__nor2_1 _08554_ (.A(\core.CPU_dmem_rd_data_a5[31] ),
    .B(net535),
    .Y(_03623_));
 sky130_fd_sc_hd__a21oi_1 _08555_ (.A1(net535),
    .A2(net476),
    .B1(_03623_),
    .Y(_03624_));
 sky130_fd_sc_hd__a21oi_1 _08556_ (.A1(_03619_),
    .A2(_03622_),
    .B1(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__or3_1 _08558_ (.A(net428),
    .B(net365),
    .C(net364),
    .X(_03627_));
 sky130_fd_sc_hd__nand2_1 _08559_ (.A(\core.CPU_Xreg_value_a4[10][31] ),
    .B(net428),
    .Y(_03628_));
 sky130_fd_sc_hd__a21oi_1 _08560_ (.A1(_03627_),
    .A2(_03628_),
    .B1(net607),
    .Y(_00776_));
 sky130_fd_sc_hd__nor2_1 _08561_ (.A(_00037_),
    .B(_02700_),
    .Y(_03629_));
 sky130_fd_sc_hd__o21bai_1 _08562_ (.A1(_00040_),
    .A2(_03629_),
    .B1_N(_00041_),
    .Y(_03630_));
 sky130_fd_sc_hd__xnor2_1 _08563_ (.A(_00046_),
    .B(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand2b_1 _08564_ (.A_N(_00036_),
    .B(_02687_),
    .Y(_03632_));
 sky130_fd_sc_hd__a21oi_1 _08565_ (.A1(_00040_),
    .A2(_03632_),
    .B1(_00039_),
    .Y(_03633_));
 sky130_fd_sc_hd__xor2_1 _08566_ (.A(_00046_),
    .B(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__a21o_1 _08567_ (.A1(_00000_),
    .A2(_00033_),
    .B1(_00032_),
    .X(_03635_));
 sky130_fd_sc_hd__nand2_1 _08568_ (.A(\core.CPU_src1_value_a3[2] ),
    .B(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__xnor2_1 _08569_ (.A(_00043_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__a221oi_1 _08570_ (.A1(_02530_),
    .A2(_02670_),
    .B1(_03637_),
    .B2(net546),
    .C1(net609),
    .Y(_03638_));
 sky130_fd_sc_hd__a211oi_1 _08571_ (.A1(net609),
    .A2(_03634_),
    .B1(_03638_),
    .C1(net612),
    .Y(_03639_));
 sky130_fd_sc_hd__a21oi_1 _08572_ (.A1(net612),
    .A2(_03631_),
    .B1(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__nand2_1 _08573_ (.A(net611),
    .B(_03637_),
    .Y(_03641_));
 sky130_fd_sc_hd__o21ai_1 _08574_ (.A1(net611),
    .A2(_03640_),
    .B1(_03641_),
    .Y(\core.CPU_result_a3[3] ));
 sky130_fd_sc_hd__mux2i_1 _08575_ (.A0(\core.CPU_dmem_rd_data_a5[3] ),
    .A1(net372),
    .S(net535),
    .Y(_03642_));
 sky130_fd_sc_hd__nand2_1 _08576_ (.A(\core.CPU_Xreg_value_a4[10][3] ),
    .B(net428),
    .Y(_03643_));
 sky130_fd_sc_hd__o211ai_1 _08578_ (.A1(net428),
    .A2(net363),
    .B1(_03643_),
    .C1(net549),
    .Y(_00777_));
 sky130_fd_sc_hd__nand2_1 _08579_ (.A(_02667_),
    .B(net478),
    .Y(_03645_));
 sky130_fd_sc_hd__xnor2_1 _08580_ (.A(_00049_),
    .B(_02631_),
    .Y(_03646_));
 sky130_fd_sc_hd__nand2_1 _08581_ (.A(net546),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__o211ai_1 _08582_ (.A1(_03645_),
    .A2(_02748_),
    .B1(_03647_),
    .C1(net556),
    .Y(_03648_));
 sky130_fd_sc_hd__o21a_1 _08583_ (.A1(_00039_),
    .A2(_02611_),
    .B1(_00046_),
    .X(_03649_));
 sky130_fd_sc_hd__nor3_1 _08584_ (.A(_00052_),
    .B(_00045_),
    .C(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__o21ai_0 _08585_ (.A1(_02613_),
    .A2(_03650_),
    .B1(net609),
    .Y(_03651_));
 sky130_fd_sc_hd__a21oi_1 _08586_ (.A1(_03648_),
    .A2(_03651_),
    .B1(net612),
    .Y(_03652_));
 sky130_fd_sc_hd__nor2_1 _08587_ (.A(_00041_),
    .B(_02594_),
    .Y(_03653_));
 sky130_fd_sc_hd__nor2_1 _08588_ (.A(_00046_),
    .B(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__nor3_1 _08589_ (.A(_00047_),
    .B(_00052_),
    .C(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__o21ai_0 _08590_ (.A1(_00047_),
    .A2(_03654_),
    .B1(_00052_),
    .Y(_03656_));
 sky130_fd_sc_hd__nor3b_1 _08591_ (.A(_03655_),
    .B(net555),
    .C_N(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__nand2_1 _08592_ (.A(net611),
    .B(_03646_),
    .Y(_03658_));
 sky130_fd_sc_hd__o31a_1 _08593_ (.A1(net611),
    .A2(_03652_),
    .A3(_03657_),
    .B1(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__nand2_1 _08594_ (.A(net536),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__o21ai_2 _08595_ (.A1(\core.CPU_dmem_rd_data_a5[4] ),
    .A2(net536),
    .B1(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__or2_0 _08596_ (.A(net607),
    .B(net352),
    .X(_03662_));
 sky130_fd_sc_hd__nand3_1 _08597_ (.A(\core.CPU_Xreg_value_a4[10][4] ),
    .B(net549),
    .C(net428),
    .Y(_03663_));
 sky130_fd_sc_hd__o21ai_0 _08598_ (.A1(net428),
    .A2(_03662_),
    .B1(_03663_),
    .Y(_00778_));
 sky130_fd_sc_hd__inv_1 _08599_ (.A(_00056_),
    .Y(_03664_));
 sky130_fd_sc_hd__nor2_1 _08600_ (.A(_02690_),
    .B(_02779_),
    .Y(_03665_));
 sky130_fd_sc_hd__xnor2_1 _08601_ (.A(_03664_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__a21oi_1 _08602_ (.A1(net609),
    .A2(_03666_),
    .B1(_02853_),
    .Y(_03667_));
 sky130_fd_sc_hd__nor2_1 _08603_ (.A(_02654_),
    .B(_02655_),
    .Y(_03668_));
 sky130_fd_sc_hd__a21oi_1 _08604_ (.A1(_00049_),
    .A2(_03668_),
    .B1(_00048_),
    .Y(_03669_));
 sky130_fd_sc_hd__xor2_1 _08605_ (.A(_00059_),
    .B(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__o221ai_1 _08606_ (.A1(_03645_),
    .A2(_02801_),
    .B1(_03670_),
    .B2(_02540_),
    .C1(net556),
    .Y(_03671_));
 sky130_fd_sc_hd__nand2_1 _08607_ (.A(_02704_),
    .B(_03178_),
    .Y(_03672_));
 sky130_fd_sc_hd__xnor2_1 _08608_ (.A(_03664_),
    .B(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__o22ai_1 _08609_ (.A1(_02804_),
    .A2(_03673_),
    .B1(_03670_),
    .B2(net557),
    .Y(_03674_));
 sky130_fd_sc_hd__a21oi_1 _08610_ (.A1(_03667_),
    .A2(_03671_),
    .B1(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__nand2_1 _08611_ (.A(\core.CPU_dmem_rd_data_a5[5] ),
    .B(net562),
    .Y(_03676_));
 sky130_fd_sc_hd__o21ai_1 _08612_ (.A1(net562),
    .A2(_03675_),
    .B1(_03676_),
    .Y(_03677_));
 sky130_fd_sc_hd__nand2_1 _08613_ (.A(_02558_),
    .B(net371),
    .Y(_03678_));
 sky130_fd_sc_hd__nand2_1 _08614_ (.A(\core.CPU_Xreg_value_a4[10][5] ),
    .B(net428),
    .Y(_03679_));
 sky130_fd_sc_hd__a21oi_1 _08615_ (.A1(_03678_),
    .A2(_03679_),
    .B1(net607),
    .Y(_00779_));
 sky130_fd_sc_hd__a22o_1 _08616_ (.A1(_02629_),
    .A2(_02630_),
    .B1(_02631_),
    .B2(_02632_),
    .X(_03680_));
 sky130_fd_sc_hd__xor2_1 _08617_ (.A(_00067_),
    .B(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__o21ai_0 _08618_ (.A1(_02540_),
    .A2(_03681_),
    .B1(net556),
    .Y(_03682_));
 sky130_fd_sc_hd__a31oi_1 _08619_ (.A1(_02667_),
    .A2(net478),
    .A3(_02838_),
    .B1(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__o21ai_0 _08620_ (.A1(_00051_),
    .A2(_02613_),
    .B1(_00056_),
    .Y(_03684_));
 sky130_fd_sc_hd__nor2_1 _08621_ (.A(_00062_),
    .B(_00055_),
    .Y(_03685_));
 sky130_fd_sc_hd__a21oi_1 _08622_ (.A1(_03684_),
    .A2(_03685_),
    .B1(_02843_),
    .Y(_03686_));
 sky130_fd_sc_hd__o21ai_0 _08623_ (.A1(net556),
    .A2(_03686_),
    .B1(net555),
    .Y(_03687_));
 sky130_fd_sc_hd__o211ai_1 _08624_ (.A1(_02594_),
    .A2(_02595_),
    .B1(_02596_),
    .C1(_02597_),
    .Y(_03688_));
 sky130_fd_sc_hd__a21oi_1 _08625_ (.A1(_00053_),
    .A2(_03664_),
    .B1(_00057_),
    .Y(_03689_));
 sky130_fd_sc_hd__nand2_1 _08626_ (.A(_03688_),
    .B(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__xnor2_1 _08627_ (.A(_02707_),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__o22ai_1 _08628_ (.A1(_03683_),
    .A2(_03687_),
    .B1(_03691_),
    .B2(net555),
    .Y(_03692_));
 sky130_fd_sc_hd__nor2_1 _08629_ (.A(net557),
    .B(_03681_),
    .Y(_03693_));
 sky130_fd_sc_hd__a21oi_1 _08630_ (.A1(net557),
    .A2(_03692_),
    .B1(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__nand2_1 _08631_ (.A(net536),
    .B(_03694_),
    .Y(_03695_));
 sky130_fd_sc_hd__o211ai_1 _08632_ (.A1(\core.CPU_dmem_rd_data_a5[6] ),
    .A2(net536),
    .B1(_03695_),
    .C1(_02644_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand3_1 _08634_ (.A(\core.CPU_Xreg_value_a4[10][6] ),
    .B(_02644_),
    .C(_02563_),
    .Y(_03698_));
 sky130_fd_sc_hd__o21ai_0 _08635_ (.A1(_02563_),
    .A2(net344),
    .B1(_03698_),
    .Y(_00780_));
 sky130_fd_sc_hd__xor2_1 _08636_ (.A(_00070_),
    .B(_02710_),
    .X(_03699_));
 sky130_fd_sc_hd__xor2_1 _08637_ (.A(_00065_),
    .B(_02770_),
    .X(_03700_));
 sky130_fd_sc_hd__o21ai_0 _08638_ (.A1(_02614_),
    .A2(_03665_),
    .B1(_02691_),
    .Y(_03701_));
 sky130_fd_sc_hd__xor2_1 _08639_ (.A(_00070_),
    .B(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__o21ai_0 _08640_ (.A1(_03087_),
    .A2(_03700_),
    .B1(net547),
    .Y(_03703_));
 sky130_fd_sc_hd__nor3_1 _08641_ (.A(net609),
    .B(_03645_),
    .C(_02894_),
    .Y(_03704_));
 sky130_fd_sc_hd__a211oi_1 _08642_ (.A1(net609),
    .A2(_03702_),
    .B1(_03703_),
    .C1(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__a221oi_1 _08643_ (.A1(net476),
    .A2(_03699_),
    .B1(_03700_),
    .B2(net611),
    .C1(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__mux2i_1 _08644_ (.A0(\core.CPU_dmem_rd_data_a5[7] ),
    .A1(_03706_),
    .S(net536),
    .Y(_03707_));
 sky130_fd_sc_hd__o21ai_0 _08645_ (.A1(\core.CPU_Xreg_value_a4[10][7] ),
    .A2(net429),
    .B1(net552),
    .Y(_03708_));
 sky130_fd_sc_hd__a21oi_1 _08646_ (.A1(net429),
    .A2(net362),
    .B1(_03708_),
    .Y(_00781_));
 sky130_fd_sc_hd__xor2_1 _08647_ (.A(_00073_),
    .B(_02635_),
    .X(_03709_));
 sky130_fd_sc_hd__a22oi_1 _08648_ (.A1(_03286_),
    .A2(_03423_),
    .B1(_03709_),
    .B2(net546),
    .Y(_03710_));
 sky130_fd_sc_hd__nor2_1 _08649_ (.A(_02539_),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__nand2_1 _08650_ (.A(_02601_),
    .B(_02602_),
    .Y(_03712_));
 sky130_fd_sc_hd__a211oi_1 _08651_ (.A1(_03688_),
    .A2(_03689_),
    .B1(_00062_),
    .C1(_00070_),
    .Y(_03713_));
 sky130_fd_sc_hd__o21a_1 _08652_ (.A1(_03712_),
    .A2(_03713_),
    .B1(_00076_),
    .X(_03714_));
 sky130_fd_sc_hd__nor3_1 _08653_ (.A(_00076_),
    .B(_03712_),
    .C(_03713_),
    .Y(_03715_));
 sky130_fd_sc_hd__o21ai_0 _08654_ (.A1(_03714_),
    .A2(_03715_),
    .B1(net612),
    .Y(_03716_));
 sky130_fd_sc_hd__inv_1 _08655_ (.A(_00069_),
    .Y(_03717_));
 sky130_fd_sc_hd__o21ai_0 _08656_ (.A1(_00061_),
    .A2(_02843_),
    .B1(_00070_),
    .Y(_03718_));
 sky130_fd_sc_hd__a211o_1 _08657_ (.A1(_03717_),
    .A2(_03718_),
    .B1(_02609_),
    .C1(_00076_),
    .X(_03719_));
 sky130_fd_sc_hd__nand4_1 _08658_ (.A(_00076_),
    .B(_03717_),
    .C(_02681_),
    .D(_03718_),
    .Y(_03720_));
 sky130_fd_sc_hd__nor2_1 _08659_ (.A(net557),
    .B(_03709_),
    .Y(_03721_));
 sky130_fd_sc_hd__a41oi_1 _08660_ (.A1(net557),
    .A2(_03716_),
    .A3(_03719_),
    .A4(_03720_),
    .B1(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__nor3_1 _08661_ (.A(net562),
    .B(_03711_),
    .C(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__nor2_1 _08662_ (.A(\core.CPU_dmem_rd_data_a5[8] ),
    .B(net536),
    .Y(_03724_));
 sky130_fd_sc_hd__nor3_2 _08663_ (.A(\core.CPU_reset_a3 ),
    .B(_03723_),
    .C(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__nand2_1 _08664_ (.A(net429),
    .B(net351),
    .Y(_03726_));
 sky130_fd_sc_hd__nand3_1 _08666_ (.A(\core.CPU_Xreg_value_a4[10][8] ),
    .B(net551),
    .C(_02563_),
    .Y(_03728_));
 sky130_fd_sc_hd__nand2_1 _08667_ (.A(_03726_),
    .B(_03728_),
    .Y(_00782_));
 sky130_fd_sc_hd__o21a_1 _08668_ (.A1(_02781_),
    .A2(_02785_),
    .B1(_00080_),
    .X(_03729_));
 sky130_fd_sc_hd__nor3_1 _08669_ (.A(_00080_),
    .B(_02781_),
    .C(_02785_),
    .Y(_03730_));
 sky130_fd_sc_hd__o21ai_0 _08670_ (.A1(_03729_),
    .A2(_03730_),
    .B1(_02681_),
    .Y(_03731_));
 sky130_fd_sc_hd__or3_1 _08671_ (.A(_00080_),
    .B(_03180_),
    .C(_03182_),
    .X(_03732_));
 sky130_fd_sc_hd__o21ai_0 _08672_ (.A1(_03180_),
    .A2(_03182_),
    .B1(_00080_),
    .Y(_03733_));
 sky130_fd_sc_hd__nand3_1 _08673_ (.A(net612),
    .B(_03732_),
    .C(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _08674_ (.A(_03731_),
    .B(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand3_1 _08675_ (.A(net548),
    .B(_02588_),
    .C(_02799_),
    .Y(_03736_));
 sky130_fd_sc_hd__o21ai_0 _08676_ (.A1(net480),
    .A2(_02989_),
    .B1(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__a21oi_1 _08677_ (.A1(_02667_),
    .A2(_03737_),
    .B1(_02539_),
    .Y(_03738_));
 sky130_fd_sc_hd__xnor2_1 _08678_ (.A(_00083_),
    .B(_02771_),
    .Y(_03739_));
 sky130_fd_sc_hd__a31oi_1 _08679_ (.A1(net546),
    .A2(_03731_),
    .A3(_03734_),
    .B1(net611),
    .Y(_03740_));
 sky130_fd_sc_hd__o32ai_1 _08680_ (.A1(net611),
    .A2(_03735_),
    .A3(_03738_),
    .B1(_03739_),
    .B2(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__nor2_1 _08681_ (.A(net562),
    .B(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__nor2_1 _08682_ (.A(\core.CPU_dmem_rd_data_a5[9] ),
    .B(net536),
    .Y(_03743_));
 sky130_fd_sc_hd__or3_1 _08683_ (.A(\core.CPU_reset_a3 ),
    .B(_03742_),
    .C(_03743_),
    .X(_03744_));
 sky130_fd_sc_hd__nand3_1 _08685_ (.A(\core.CPU_Xreg_value_a4[10][9] ),
    .B(net552),
    .C(net428),
    .Y(_03746_));
 sky130_fd_sc_hd__o21ai_0 _08686_ (.A1(net428),
    .A2(_03744_),
    .B1(_03746_),
    .Y(_00783_));
 sky130_fd_sc_hd__a21o_1 _08687_ (.A1(net535),
    .A2(net394),
    .B1(net440),
    .X(_03747_));
 sky130_fd_sc_hd__and3_1 _08688_ (.A(\core.CPU_rd_a3[0] ),
    .B(\core.CPU_rd_a3[1] ),
    .C(net535),
    .X(_03748_));
 sky130_fd_sc_hd__and3_1 _08689_ (.A(\core.CPU_rd_a5[0] ),
    .B(\core.CPU_rd_a5[1] ),
    .C(_01114_),
    .X(_03749_));
 sky130_fd_sc_hd__o21a_1 _08690_ (.A1(_03748_),
    .A2(_03749_),
    .B1(_02556_),
    .X(_03750_));
 sky130_fd_sc_hd__nand2_2 _08691_ (.A(_02561_),
    .B(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__nand2_1 _08695_ (.A(\core.CPU_Xreg_value_a4[11][0] ),
    .B(_03751_),
    .Y(_03755_));
 sky130_fd_sc_hd__o211ai_1 _08696_ (.A1(_03747_),
    .A2(_03751_),
    .B1(_03755_),
    .C1(net549),
    .Y(_00784_));
 sky130_fd_sc_hd__nand3_1 _08698_ (.A(\core.CPU_Xreg_value_a4[11][10] ),
    .B(net550),
    .C(_03751_),
    .Y(_03757_));
 sky130_fd_sc_hd__o21ai_0 _08699_ (.A1(net348),
    .A2(_03751_),
    .B1(_03757_),
    .Y(_00785_));
 sky130_fd_sc_hd__nand3_1 _08700_ (.A(\core.CPU_Xreg_value_a4[11][11] ),
    .B(net550),
    .C(_03751_),
    .Y(_03758_));
 sky130_fd_sc_hd__o21ai_0 _08701_ (.A1(net361),
    .A2(_03751_),
    .B1(_03758_),
    .Y(_00786_));
 sky130_fd_sc_hd__o21ai_0 _08703_ (.A1(_03748_),
    .A2(_03749_),
    .B1(_02556_),
    .Y(_03760_));
 sky130_fd_sc_hd__nor2_2 _08704_ (.A(_02550_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__nand2_1 _08706_ (.A(net360),
    .B(net425),
    .Y(_03763_));
 sky130_fd_sc_hd__nand2_1 _08707_ (.A(\core.CPU_Xreg_value_a4[11][12] ),
    .B(net426),
    .Y(_03764_));
 sky130_fd_sc_hd__a21oi_1 _08708_ (.A1(_03763_),
    .A2(_03764_),
    .B1(net606),
    .Y(_00787_));
 sky130_fd_sc_hd__nand3_1 _08709_ (.A(\core.CPU_Xreg_value_a4[11][13] ),
    .B(net552),
    .C(net426),
    .Y(_03765_));
 sky130_fd_sc_hd__o31ai_1 _08710_ (.A1(_02811_),
    .A2(net439),
    .A3(net426),
    .B1(_03765_),
    .Y(_00788_));
 sky130_fd_sc_hd__nand3_1 _08711_ (.A(\core.CPU_Xreg_value_a4[11][14] ),
    .B(net549),
    .C(_03751_),
    .Y(_03766_));
 sky130_fd_sc_hd__o21ai_0 _08712_ (.A1(net347),
    .A2(_03751_),
    .B1(_03766_),
    .Y(_00789_));
 sky130_fd_sc_hd__nand3_1 _08714_ (.A(\core.CPU_Xreg_value_a4[11][15] ),
    .B(net551),
    .C(net426),
    .Y(_03768_));
 sky130_fd_sc_hd__o21ai_0 _08715_ (.A1(_02911_),
    .A2(net426),
    .B1(_03768_),
    .Y(_00790_));
 sky130_fd_sc_hd__o21ai_0 _08718_ (.A1(\core.CPU_Xreg_value_a4[11][16] ),
    .A2(net425),
    .B1(net551),
    .Y(_03771_));
 sky130_fd_sc_hd__a21oi_1 _08719_ (.A1(net346),
    .A2(net425),
    .B1(_03771_),
    .Y(_00791_));
 sky130_fd_sc_hd__nand2_1 _08721_ (.A(_02961_),
    .B(net425),
    .Y(_03773_));
 sky130_fd_sc_hd__nand3_1 _08722_ (.A(\core.CPU_Xreg_value_a4[11][17] ),
    .B(net552),
    .C(net426),
    .Y(_03774_));
 sky130_fd_sc_hd__o221ai_1 _08723_ (.A1(_03006_),
    .A2(net426),
    .B1(_03773_),
    .B2(_03003_),
    .C1(_03774_),
    .Y(_00792_));
 sky130_fd_sc_hd__nand3_1 _08726_ (.A(\core.CPU_Xreg_value_a4[11][18] ),
    .B(net552),
    .C(net426),
    .Y(_03777_));
 sky130_fd_sc_hd__o221ai_1 _08727_ (.A1(_03043_),
    .A2(net426),
    .B1(_03773_),
    .B2(net359),
    .C1(_03777_),
    .Y(_00793_));
 sky130_fd_sc_hd__o21ai_0 _08729_ (.A1(\core.CPU_Xreg_value_a4[11][19] ),
    .A2(net425),
    .B1(_02644_),
    .Y(_03779_));
 sky130_fd_sc_hd__a21oi_1 _08730_ (.A1(net358),
    .A2(net425),
    .B1(_03779_),
    .Y(_00794_));
 sky130_fd_sc_hd__nor3_1 _08732_ (.A(\core.CPU_Xreg_value_a4[11][1] ),
    .B(net607),
    .C(_03761_),
    .Y(_03781_));
 sky130_fd_sc_hd__a31oi_1 _08733_ (.A1(_02644_),
    .A2(net375),
    .A3(_03761_),
    .B1(_03781_),
    .Y(_00795_));
 sky130_fd_sc_hd__nand3_1 _08734_ (.A(\core.CPU_Xreg_value_a4[11][20] ),
    .B(net549),
    .C(_03751_),
    .Y(_03782_));
 sky130_fd_sc_hd__o21ai_0 _08735_ (.A1(net357),
    .A2(_03751_),
    .B1(_03782_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand3_1 _08736_ (.A(\core.CPU_Xreg_value_a4[11][21] ),
    .B(net550),
    .C(_03751_),
    .Y(_03783_));
 sky130_fd_sc_hd__o21ai_0 _08737_ (.A1(net356),
    .A2(_03751_),
    .B1(_03783_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_1 _08738_ (.A(\core.CPU_Xreg_value_a4[11][22] ),
    .B(net426),
    .Y(_03784_));
 sky130_fd_sc_hd__nand2_1 _08740_ (.A(net355),
    .B(net425),
    .Y(_03786_));
 sky130_fd_sc_hd__a21oi_1 _08741_ (.A1(_03784_),
    .A2(_03786_),
    .B1(net607),
    .Y(_00798_));
 sky130_fd_sc_hd__nand2_1 _08743_ (.A(net368),
    .B(net425),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_1 _08744_ (.A(\core.CPU_Xreg_value_a4[11][23] ),
    .B(net426),
    .Y(_03789_));
 sky130_fd_sc_hd__a21oi_1 _08745_ (.A1(_03788_),
    .A2(_03789_),
    .B1(net606),
    .Y(_00799_));
 sky130_fd_sc_hd__o21ai_0 _08747_ (.A1(\core.CPU_Xreg_value_a4[11][24] ),
    .A2(net425),
    .B1(net552),
    .Y(_03791_));
 sky130_fd_sc_hd__a21oi_2 _08748_ (.A1(_03309_),
    .A2(net425),
    .B1(_03791_),
    .Y(_00800_));
 sky130_fd_sc_hd__o21ai_0 _08750_ (.A1(\core.CPU_Xreg_value_a4[11][25] ),
    .A2(net425),
    .B1(_02644_),
    .Y(_03793_));
 sky130_fd_sc_hd__a21oi_1 _08751_ (.A1(net354),
    .A2(net425),
    .B1(_03793_),
    .Y(_00801_));
 sky130_fd_sc_hd__o21ai_0 _08753_ (.A1(\core.CPU_Xreg_value_a4[11][26] ),
    .A2(net425),
    .B1(net551),
    .Y(_03795_));
 sky130_fd_sc_hd__a21oi_1 _08754_ (.A1(_03389_),
    .A2(net425),
    .B1(_03795_),
    .Y(_00802_));
 sky130_fd_sc_hd__nor2_1 _08755_ (.A(_01114_),
    .B(net426),
    .Y(_03796_));
 sky130_fd_sc_hd__nand2_1 _08757_ (.A(net436),
    .B(net425),
    .Y(_03798_));
 sky130_fd_sc_hd__o21ai_0 _08758_ (.A1(\core.CPU_Xreg_value_a4[11][27] ),
    .A2(net425),
    .B1(_03798_),
    .Y(_03799_));
 sky130_fd_sc_hd__a311oi_1 _08759_ (.A1(net353),
    .A2(_03431_),
    .A3(_03796_),
    .B1(_03799_),
    .C1(net606),
    .Y(_00803_));
 sky130_fd_sc_hd__nand3_1 _08762_ (.A(_03474_),
    .B(_03475_),
    .C(net425),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_1 _08763_ (.A(\core.CPU_Xreg_value_a4[11][28] ),
    .B(net426),
    .Y(_03803_));
 sky130_fd_sc_hd__a21oi_1 _08765_ (.A1(_03802_),
    .A2(_03803_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_00804_));
 sky130_fd_sc_hd__nand3_1 _08766_ (.A(\core.CPU_Xreg_value_a4[11][29] ),
    .B(net549),
    .C(_03751_),
    .Y(_03805_));
 sky130_fd_sc_hd__o21ai_0 _08767_ (.A1(_03523_),
    .A2(_03751_),
    .B1(_03805_),
    .Y(_00805_));
 sky130_fd_sc_hd__nor2_1 _08768_ (.A(net373),
    .B(_03751_),
    .Y(_03806_));
 sky130_fd_sc_hd__o21ai_0 _08769_ (.A1(\core.CPU_Xreg_value_a4[11][2] ),
    .A2(_03761_),
    .B1(_02644_),
    .Y(_03807_));
 sky130_fd_sc_hd__nor2_1 _08770_ (.A(_03806_),
    .B(_03807_),
    .Y(_00806_));
 sky130_fd_sc_hd__o21ai_0 _08773_ (.A1(\core.CPU_Xreg_value_a4[11][30] ),
    .A2(net425),
    .B1(_02644_),
    .Y(_03810_));
 sky130_fd_sc_hd__a21oi_1 _08774_ (.A1(net345),
    .A2(net425),
    .B1(_03810_),
    .Y(_00807_));
 sky130_fd_sc_hd__or3_1 _08775_ (.A(net365),
    .B(net364),
    .C(_03751_),
    .X(_03811_));
 sky130_fd_sc_hd__nand2_1 _08776_ (.A(\core.CPU_Xreg_value_a4[11][31] ),
    .B(_03751_),
    .Y(_03812_));
 sky130_fd_sc_hd__a21oi_1 _08777_ (.A1(_03811_),
    .A2(_03812_),
    .B1(net607),
    .Y(_00808_));
 sky130_fd_sc_hd__nand2_1 _08778_ (.A(\core.CPU_Xreg_value_a4[11][3] ),
    .B(_03751_),
    .Y(_03813_));
 sky130_fd_sc_hd__o211ai_1 _08779_ (.A1(net363),
    .A2(_03751_),
    .B1(_03813_),
    .C1(net549),
    .Y(_00809_));
 sky130_fd_sc_hd__nand3_1 _08780_ (.A(\core.CPU_Xreg_value_a4[11][4] ),
    .B(net549),
    .C(_03751_),
    .Y(_03814_));
 sky130_fd_sc_hd__o21ai_0 _08781_ (.A1(_03662_),
    .A2(_03751_),
    .B1(_03814_),
    .Y(_00810_));
 sky130_fd_sc_hd__nand2_1 _08783_ (.A(net371),
    .B(_03761_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2_1 _08784_ (.A(\core.CPU_Xreg_value_a4[11][5] ),
    .B(_03751_),
    .Y(_03817_));
 sky130_fd_sc_hd__a21oi_1 _08785_ (.A1(_03816_),
    .A2(_03817_),
    .B1(net607),
    .Y(_00811_));
 sky130_fd_sc_hd__nand3_1 _08786_ (.A(\core.CPU_Xreg_value_a4[11][6] ),
    .B(_02644_),
    .C(net426),
    .Y(_03818_));
 sky130_fd_sc_hd__o21ai_0 _08787_ (.A1(net344),
    .A2(net426),
    .B1(_03818_),
    .Y(_00812_));
 sky130_fd_sc_hd__o21ai_0 _08789_ (.A1(\core.CPU_Xreg_value_a4[11][7] ),
    .A2(net425),
    .B1(net552),
    .Y(_03820_));
 sky130_fd_sc_hd__a21oi_1 _08790_ (.A1(net362),
    .A2(net425),
    .B1(_03820_),
    .Y(_00813_));
 sky130_fd_sc_hd__nand2_1 _08792_ (.A(net351),
    .B(net425),
    .Y(_03822_));
 sky130_fd_sc_hd__nand3_1 _08793_ (.A(\core.CPU_Xreg_value_a4[11][8] ),
    .B(net551),
    .C(net426),
    .Y(_03823_));
 sky130_fd_sc_hd__nand2_1 _08794_ (.A(_03822_),
    .B(_03823_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand3_1 _08795_ (.A(\core.CPU_Xreg_value_a4[11][9] ),
    .B(net552),
    .C(net426),
    .Y(_03824_));
 sky130_fd_sc_hd__o21ai_0 _08796_ (.A1(_03744_),
    .A2(net426),
    .B1(_03824_),
    .Y(_00815_));
 sky130_fd_sc_hd__a31oi_1 _08797_ (.A1(\core.CPU_rd_valid_a3 ),
    .A2(_01115_),
    .A3(_02555_),
    .B1(\core.CPU_valid_load_a5 ),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2b_1 _08798_ (.A_N(\core.CPU_rd_a5[3] ),
    .B(\core.CPU_rd_a5[4] ),
    .Y(_03826_));
 sky130_fd_sc_hd__or3_1 _08799_ (.A(\core.CPU_rd_a3[3] ),
    .B(_02548_),
    .C(_01114_),
    .X(_03827_));
 sky130_fd_sc_hd__o21a_1 _08800_ (.A1(net535),
    .A2(_03826_),
    .B1(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__nor3_1 _08801_ (.A(\core.CPU_rd_a5[0] ),
    .B(\core.CPU_rd_a5[1] ),
    .C(net535),
    .Y(_03829_));
 sky130_fd_sc_hd__a21oi_1 _08802_ (.A1(net535),
    .A2(_02553_),
    .B1(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__nor3_2 _08803_ (.A(_03825_),
    .B(_03828_),
    .C(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand2_1 _08805_ (.A(_02545_),
    .B(net424),
    .Y(_03833_));
 sky130_fd_sc_hd__o21ai_0 _08806_ (.A1(net535),
    .A2(_03826_),
    .B1(_03827_),
    .Y(_03834_));
 sky130_fd_sc_hd__nor2_1 _08807_ (.A(_03825_),
    .B(_03830_),
    .Y(_03835_));
 sky130_fd_sc_hd__nand2_2 _08808_ (.A(_03834_),
    .B(_03835_),
    .Y(_03836_));
 sky130_fd_sc_hd__nand2_1 _08811_ (.A(\core.CPU_Xreg_value_a4[16][0] ),
    .B(net390),
    .Y(_03839_));
 sky130_fd_sc_hd__a21oi_1 _08812_ (.A1(_03833_),
    .A2(_03839_),
    .B1(net607),
    .Y(_00816_));
 sky130_fd_sc_hd__nand3_1 _08815_ (.A(\core.CPU_Xreg_value_a4[16][10] ),
    .B(net550),
    .C(net390),
    .Y(_03842_));
 sky130_fd_sc_hd__o21ai_0 _08816_ (.A1(net348),
    .A2(net390),
    .B1(_03842_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand3_1 _08817_ (.A(\core.CPU_Xreg_value_a4[16][11] ),
    .B(net550),
    .C(net390),
    .Y(_03843_));
 sky130_fd_sc_hd__o21ai_0 _08818_ (.A1(net361),
    .A2(net390),
    .B1(_03843_),
    .Y(_00818_));
 sky130_fd_sc_hd__nand2_1 _08820_ (.A(net360),
    .B(net424),
    .Y(_03845_));
 sky130_fd_sc_hd__nand2_1 _08821_ (.A(\core.CPU_Xreg_value_a4[16][12] ),
    .B(_03836_),
    .Y(_03846_));
 sky130_fd_sc_hd__a21oi_1 _08822_ (.A1(_03845_),
    .A2(_03846_),
    .B1(net606),
    .Y(_00819_));
 sky130_fd_sc_hd__nand3_1 _08823_ (.A(\core.CPU_Xreg_value_a4[16][13] ),
    .B(net552),
    .C(_03836_),
    .Y(_03847_));
 sky130_fd_sc_hd__o31ai_1 _08824_ (.A1(_02811_),
    .A2(net439),
    .A3(_03836_),
    .B1(_03847_),
    .Y(_00820_));
 sky130_fd_sc_hd__nand3_1 _08825_ (.A(\core.CPU_Xreg_value_a4[16][14] ),
    .B(net549),
    .C(net390),
    .Y(_03848_));
 sky130_fd_sc_hd__o21ai_0 _08826_ (.A1(net347),
    .A2(net390),
    .B1(_03848_),
    .Y(_00821_));
 sky130_fd_sc_hd__nand3_1 _08828_ (.A(\core.CPU_Xreg_value_a4[16][15] ),
    .B(net551),
    .C(_03836_),
    .Y(_03850_));
 sky130_fd_sc_hd__o21ai_0 _08829_ (.A1(_02911_),
    .A2(_03836_),
    .B1(_03850_),
    .Y(_00822_));
 sky130_fd_sc_hd__o21ai_0 _08830_ (.A1(\core.CPU_Xreg_value_a4[16][16] ),
    .A2(net424),
    .B1(net551),
    .Y(_03851_));
 sky130_fd_sc_hd__a21oi_1 _08831_ (.A1(net346),
    .A2(net424),
    .B1(_03851_),
    .Y(_00823_));
 sky130_fd_sc_hd__nand2_1 _08832_ (.A(_02961_),
    .B(net424),
    .Y(_03852_));
 sky130_fd_sc_hd__nand3_1 _08833_ (.A(\core.CPU_Xreg_value_a4[16][17] ),
    .B(net552),
    .C(_03836_),
    .Y(_03853_));
 sky130_fd_sc_hd__o221ai_1 _08834_ (.A1(_03006_),
    .A2(_03836_),
    .B1(_03852_),
    .B2(_03003_),
    .C1(_03853_),
    .Y(_00824_));
 sky130_fd_sc_hd__nand3_1 _08835_ (.A(\core.CPU_Xreg_value_a4[16][18] ),
    .B(net552),
    .C(_03836_),
    .Y(_03854_));
 sky130_fd_sc_hd__o221ai_1 _08836_ (.A1(_03043_),
    .A2(_03836_),
    .B1(_03852_),
    .B2(net359),
    .C1(_03854_),
    .Y(_00825_));
 sky130_fd_sc_hd__o21ai_0 _08837_ (.A1(\core.CPU_Xreg_value_a4[16][19] ),
    .A2(net424),
    .B1(_02644_),
    .Y(_03855_));
 sky130_fd_sc_hd__a21oi_1 _08838_ (.A1(net358),
    .A2(net424),
    .B1(_03855_),
    .Y(_00826_));
 sky130_fd_sc_hd__o21ai_0 _08839_ (.A1(\core.CPU_Xreg_value_a4[16][1] ),
    .A2(net424),
    .B1(_02644_),
    .Y(_03856_));
 sky130_fd_sc_hd__a21oi_1 _08840_ (.A1(net375),
    .A2(net424),
    .B1(_03856_),
    .Y(_00827_));
 sky130_fd_sc_hd__nand3_1 _08841_ (.A(\core.CPU_Xreg_value_a4[16][20] ),
    .B(net549),
    .C(net390),
    .Y(_03857_));
 sky130_fd_sc_hd__o21ai_0 _08842_ (.A1(net357),
    .A2(net390),
    .B1(_03857_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand3_1 _08843_ (.A(\core.CPU_Xreg_value_a4[16][21] ),
    .B(net550),
    .C(net390),
    .Y(_03858_));
 sky130_fd_sc_hd__o21ai_0 _08844_ (.A1(net356),
    .A2(net390),
    .B1(_03858_),
    .Y(_00829_));
 sky130_fd_sc_hd__nand2_1 _08845_ (.A(\core.CPU_Xreg_value_a4[16][22] ),
    .B(net390),
    .Y(_03859_));
 sky130_fd_sc_hd__nand2_1 _08846_ (.A(net355),
    .B(net424),
    .Y(_03860_));
 sky130_fd_sc_hd__a21oi_1 _08847_ (.A1(_03859_),
    .A2(_03860_),
    .B1(net607),
    .Y(_00830_));
 sky130_fd_sc_hd__nand2_1 _08848_ (.A(net368),
    .B(net424),
    .Y(_03861_));
 sky130_fd_sc_hd__nand2_1 _08849_ (.A(\core.CPU_Xreg_value_a4[16][23] ),
    .B(_03836_),
    .Y(_03862_));
 sky130_fd_sc_hd__a21oi_1 _08850_ (.A1(_03861_),
    .A2(_03862_),
    .B1(net606),
    .Y(_00831_));
 sky130_fd_sc_hd__o21ai_0 _08851_ (.A1(\core.CPU_Xreg_value_a4[16][24] ),
    .A2(net424),
    .B1(net552),
    .Y(_03863_));
 sky130_fd_sc_hd__a21oi_2 _08852_ (.A1(_03309_),
    .A2(net424),
    .B1(_03863_),
    .Y(_00832_));
 sky130_fd_sc_hd__o21ai_0 _08853_ (.A1(\core.CPU_Xreg_value_a4[16][25] ),
    .A2(net424),
    .B1(_02644_),
    .Y(_03864_));
 sky130_fd_sc_hd__a21oi_1 _08854_ (.A1(net354),
    .A2(net424),
    .B1(_03864_),
    .Y(_00833_));
 sky130_fd_sc_hd__o21ai_0 _08855_ (.A1(\core.CPU_Xreg_value_a4[16][26] ),
    .A2(net424),
    .B1(net551),
    .Y(_03865_));
 sky130_fd_sc_hd__a21oi_1 _08856_ (.A1(_03389_),
    .A2(net424),
    .B1(_03865_),
    .Y(_00834_));
 sky130_fd_sc_hd__nor2_1 _08857_ (.A(_01114_),
    .B(_03836_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _08858_ (.A(net436),
    .B(net424),
    .Y(_03867_));
 sky130_fd_sc_hd__o21ai_0 _08859_ (.A1(\core.CPU_Xreg_value_a4[16][27] ),
    .A2(net424),
    .B1(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__a311oi_1 _08860_ (.A1(net353),
    .A2(_03431_),
    .A3(_03866_),
    .B1(_03868_),
    .C1(net606),
    .Y(_00835_));
 sky130_fd_sc_hd__nand3_1 _08861_ (.A(_03474_),
    .B(_03475_),
    .C(net424),
    .Y(_03869_));
 sky130_fd_sc_hd__nand2_1 _08862_ (.A(\core.CPU_Xreg_value_a4[16][28] ),
    .B(_03836_),
    .Y(_03870_));
 sky130_fd_sc_hd__a21oi_1 _08863_ (.A1(_03869_),
    .A2(_03870_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_00836_));
 sky130_fd_sc_hd__nand3_1 _08864_ (.A(\core.CPU_Xreg_value_a4[16][29] ),
    .B(net549),
    .C(net390),
    .Y(_03871_));
 sky130_fd_sc_hd__o21ai_0 _08865_ (.A1(_03523_),
    .A2(net390),
    .B1(_03871_),
    .Y(_00837_));
 sky130_fd_sc_hd__nor2_1 _08866_ (.A(net373),
    .B(net390),
    .Y(_03872_));
 sky130_fd_sc_hd__o21ai_0 _08867_ (.A1(\core.CPU_Xreg_value_a4[16][2] ),
    .A2(net424),
    .B1(_02644_),
    .Y(_03873_));
 sky130_fd_sc_hd__nor2_1 _08868_ (.A(_03872_),
    .B(_03873_),
    .Y(_00838_));
 sky130_fd_sc_hd__o21ai_0 _08869_ (.A1(\core.CPU_Xreg_value_a4[16][30] ),
    .A2(net424),
    .B1(net551),
    .Y(_03874_));
 sky130_fd_sc_hd__a21oi_1 _08870_ (.A1(net345),
    .A2(net424),
    .B1(_03874_),
    .Y(_00839_));
 sky130_fd_sc_hd__or3_1 _08871_ (.A(net365),
    .B(net364),
    .C(net390),
    .X(_03875_));
 sky130_fd_sc_hd__nand2_1 _08872_ (.A(\core.CPU_Xreg_value_a4[16][31] ),
    .B(net390),
    .Y(_03876_));
 sky130_fd_sc_hd__a21oi_1 _08873_ (.A1(_03875_),
    .A2(_03876_),
    .B1(net607),
    .Y(_00840_));
 sky130_fd_sc_hd__mux2_2 _08874_ (.A0(\core.CPU_dmem_rd_data_a5[3] ),
    .A1(net372),
    .S(net535),
    .X(_03877_));
 sky130_fd_sc_hd__nand2_1 _08875_ (.A(_03877_),
    .B(net424),
    .Y(_03878_));
 sky130_fd_sc_hd__nand2_1 _08876_ (.A(\core.CPU_Xreg_value_a4[16][3] ),
    .B(net390),
    .Y(_03879_));
 sky130_fd_sc_hd__a21oi_1 _08877_ (.A1(_03878_),
    .A2(_03879_),
    .B1(net607),
    .Y(_00841_));
 sky130_fd_sc_hd__a21oi_1 _08879_ (.A1(\core.CPU_Xreg_value_a4[16][4] ),
    .A2(net390),
    .B1(net607),
    .Y(_03881_));
 sky130_fd_sc_hd__o21ai_0 _08880_ (.A1(net352),
    .A2(net390),
    .B1(_03881_),
    .Y(_00842_));
 sky130_fd_sc_hd__nand2_1 _08881_ (.A(net371),
    .B(net424),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2_1 _08882_ (.A(\core.CPU_Xreg_value_a4[16][5] ),
    .B(net390),
    .Y(_03883_));
 sky130_fd_sc_hd__a21oi_1 _08884_ (.A1(_03882_),
    .A2(_03883_),
    .B1(net607),
    .Y(_00843_));
 sky130_fd_sc_hd__nand3_1 _08885_ (.A(\core.CPU_Xreg_value_a4[16][6] ),
    .B(_02644_),
    .C(net390),
    .Y(_03885_));
 sky130_fd_sc_hd__o21ai_0 _08886_ (.A1(net344),
    .A2(net390),
    .B1(_03885_),
    .Y(_00844_));
 sky130_fd_sc_hd__o21ai_0 _08887_ (.A1(\core.CPU_Xreg_value_a4[16][7] ),
    .A2(net424),
    .B1(net551),
    .Y(_03886_));
 sky130_fd_sc_hd__a21oi_1 _08888_ (.A1(net362),
    .A2(net424),
    .B1(_03886_),
    .Y(_00845_));
 sky130_fd_sc_hd__nand2_1 _08889_ (.A(net351),
    .B(net424),
    .Y(_03887_));
 sky130_fd_sc_hd__nand3_1 _08890_ (.A(\core.CPU_Xreg_value_a4[16][8] ),
    .B(net551),
    .C(_03836_),
    .Y(_03888_));
 sky130_fd_sc_hd__nand2_1 _08891_ (.A(_03887_),
    .B(_03888_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand3_1 _08892_ (.A(\core.CPU_Xreg_value_a4[16][9] ),
    .B(net552),
    .C(_03836_),
    .Y(_03889_));
 sky130_fd_sc_hd__o21ai_0 _08893_ (.A1(_03744_),
    .A2(_03836_),
    .B1(_03889_),
    .Y(_00847_));
 sky130_fd_sc_hd__nor3b_1 _08894_ (.A(\core.CPU_rd_a3[1] ),
    .B(_01114_),
    .C_N(\core.CPU_rd_a3[0] ),
    .Y(_03890_));
 sky130_fd_sc_hd__nor3b_1 _08895_ (.A(\core.CPU_rd_a5[1] ),
    .B(net535),
    .C_N(\core.CPU_rd_a5[0] ),
    .Y(_03891_));
 sky130_fd_sc_hd__o21a_1 _08896_ (.A1(_03890_),
    .A2(_03891_),
    .B1(_02556_),
    .X(_03892_));
 sky130_fd_sc_hd__nand2_2 _08897_ (.A(_03834_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__nand2_1 _08901_ (.A(net620),
    .B(net423),
    .Y(_03897_));
 sky130_fd_sc_hd__o211ai_1 _08902_ (.A1(_03747_),
    .A2(net423),
    .B1(_03897_),
    .C1(net550),
    .Y(_00848_));
 sky130_fd_sc_hd__nand3_1 _08903_ (.A(\core.CPU_Xreg_value_a4[17][10] ),
    .B(net550),
    .C(net423),
    .Y(_03898_));
 sky130_fd_sc_hd__o21ai_0 _08904_ (.A1(net348),
    .A2(net423),
    .B1(_03898_),
    .Y(_00849_));
 sky130_fd_sc_hd__nand3_1 _08905_ (.A(\core.CPU_Xreg_value_a4[17][11] ),
    .B(net550),
    .C(net423),
    .Y(_03899_));
 sky130_fd_sc_hd__o21ai_0 _08906_ (.A1(net361),
    .A2(net423),
    .B1(_03899_),
    .Y(_00850_));
 sky130_fd_sc_hd__o21ai_0 _08907_ (.A1(_03890_),
    .A2(_03891_),
    .B1(_02556_),
    .Y(_03900_));
 sky130_fd_sc_hd__nor2_4 _08908_ (.A(_03828_),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2_1 _08910_ (.A(net360),
    .B(_03901_),
    .Y(_03903_));
 sky130_fd_sc_hd__nand2_1 _08912_ (.A(\core.CPU_Xreg_value_a4[17][12] ),
    .B(_03893_),
    .Y(_03905_));
 sky130_fd_sc_hd__a21oi_1 _08913_ (.A1(_03903_),
    .A2(_03905_),
    .B1(net607),
    .Y(_00851_));
 sky130_fd_sc_hd__nand3_1 _08915_ (.A(\core.CPU_Xreg_value_a4[17][13] ),
    .B(net552),
    .C(_03893_),
    .Y(_03907_));
 sky130_fd_sc_hd__o31ai_1 _08916_ (.A1(_02811_),
    .A2(net439),
    .A3(_03893_),
    .B1(_03907_),
    .Y(_00852_));
 sky130_fd_sc_hd__nand3_1 _08917_ (.A(\core.CPU_Xreg_value_a4[17][14] ),
    .B(net549),
    .C(net423),
    .Y(_03908_));
 sky130_fd_sc_hd__o21ai_0 _08918_ (.A1(net347),
    .A2(net423),
    .B1(_03908_),
    .Y(_00853_));
 sky130_fd_sc_hd__nand3_1 _08919_ (.A(\core.CPU_Xreg_value_a4[17][15] ),
    .B(net551),
    .C(_03893_),
    .Y(_03909_));
 sky130_fd_sc_hd__o21ai_0 _08920_ (.A1(_02911_),
    .A2(_03893_),
    .B1(_03909_),
    .Y(_00854_));
 sky130_fd_sc_hd__o21ai_0 _08923_ (.A1(\core.CPU_Xreg_value_a4[17][16] ),
    .A2(net422),
    .B1(net551),
    .Y(_03912_));
 sky130_fd_sc_hd__a21oi_1 _08924_ (.A1(net346),
    .A2(net422),
    .B1(_03912_),
    .Y(_00855_));
 sky130_fd_sc_hd__nand2_1 _08925_ (.A(_02961_),
    .B(_03901_),
    .Y(_03913_));
 sky130_fd_sc_hd__nor2_1 _08926_ (.A(_03006_),
    .B(_03893_),
    .Y(_03914_));
 sky130_fd_sc_hd__a31oi_1 _08927_ (.A1(\core.CPU_Xreg_value_a4[17][17] ),
    .A2(net552),
    .A3(_03893_),
    .B1(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__o21ai_0 _08928_ (.A1(_03003_),
    .A2(_03913_),
    .B1(_03915_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand3_1 _08929_ (.A(\core.CPU_Xreg_value_a4[17][18] ),
    .B(net552),
    .C(_03893_),
    .Y(_03916_));
 sky130_fd_sc_hd__o221ai_1 _08930_ (.A1(_03043_),
    .A2(_03893_),
    .B1(_03913_),
    .B2(net359),
    .C1(_03916_),
    .Y(_00857_));
 sky130_fd_sc_hd__o21ai_0 _08931_ (.A1(\core.CPU_Xreg_value_a4[17][19] ),
    .A2(_03901_),
    .B1(_02644_),
    .Y(_03917_));
 sky130_fd_sc_hd__a21oi_1 _08932_ (.A1(net358),
    .A2(_03901_),
    .B1(_03917_),
    .Y(_00858_));
 sky130_fd_sc_hd__o21ai_0 _08933_ (.A1(net619),
    .A2(net422),
    .B1(_02644_),
    .Y(_03918_));
 sky130_fd_sc_hd__a21oi_1 _08934_ (.A1(net375),
    .A2(net422),
    .B1(_03918_),
    .Y(_00859_));
 sky130_fd_sc_hd__nand3_1 _08936_ (.A(\core.CPU_Xreg_value_a4[17][20] ),
    .B(net549),
    .C(net423),
    .Y(_03920_));
 sky130_fd_sc_hd__o21ai_0 _08937_ (.A1(net357),
    .A2(net423),
    .B1(_03920_),
    .Y(_00860_));
 sky130_fd_sc_hd__nand3_1 _08938_ (.A(\core.CPU_Xreg_value_a4[17][21] ),
    .B(net549),
    .C(net423),
    .Y(_03921_));
 sky130_fd_sc_hd__o21ai_0 _08939_ (.A1(net356),
    .A2(net423),
    .B1(_03921_),
    .Y(_00861_));
 sky130_fd_sc_hd__nand2_1 _08940_ (.A(\core.CPU_Xreg_value_a4[17][22] ),
    .B(_03893_),
    .Y(_03922_));
 sky130_fd_sc_hd__nand2_1 _08941_ (.A(net355),
    .B(net422),
    .Y(_03923_));
 sky130_fd_sc_hd__a21oi_1 _08942_ (.A1(_03922_),
    .A2(_03923_),
    .B1(net607),
    .Y(_00862_));
 sky130_fd_sc_hd__nand2_1 _08943_ (.A(net368),
    .B(net422),
    .Y(_03924_));
 sky130_fd_sc_hd__nand2_1 _08944_ (.A(\core.CPU_Xreg_value_a4[17][23] ),
    .B(_03893_),
    .Y(_03925_));
 sky130_fd_sc_hd__a21oi_1 _08945_ (.A1(_03924_),
    .A2(_03925_),
    .B1(net606),
    .Y(_00863_));
 sky130_fd_sc_hd__o21ai_0 _08946_ (.A1(\core.CPU_Xreg_value_a4[17][24] ),
    .A2(_03901_),
    .B1(net552),
    .Y(_03926_));
 sky130_fd_sc_hd__a21oi_2 _08947_ (.A1(_03309_),
    .A2(_03901_),
    .B1(_03926_),
    .Y(_00864_));
 sky130_fd_sc_hd__nor2_1 _08948_ (.A(\core.CPU_Xreg_value_a4[17][25] ),
    .B(net422),
    .Y(_03927_));
 sky130_fd_sc_hd__a211oi_1 _08949_ (.A1(net354),
    .A2(net422),
    .B1(_03927_),
    .C1(net607),
    .Y(_00865_));
 sky130_fd_sc_hd__o21ai_0 _08950_ (.A1(\core.CPU_Xreg_value_a4[17][26] ),
    .A2(_03901_),
    .B1(net551),
    .Y(_03928_));
 sky130_fd_sc_hd__a21oi_1 _08951_ (.A1(_03389_),
    .A2(_03901_),
    .B1(_03928_),
    .Y(_00866_));
 sky130_fd_sc_hd__nor2_1 _08952_ (.A(_01114_),
    .B(_03893_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_1 _08953_ (.A(net436),
    .B(_03901_),
    .Y(_03930_));
 sky130_fd_sc_hd__o21ai_0 _08954_ (.A1(\core.CPU_Xreg_value_a4[17][27] ),
    .A2(_03901_),
    .B1(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hd__a311oi_1 _08955_ (.A1(net353),
    .A2(_03431_),
    .A3(_03929_),
    .B1(_03931_),
    .C1(net606),
    .Y(_00867_));
 sky130_fd_sc_hd__nand3_1 _08956_ (.A(_03474_),
    .B(_03475_),
    .C(_03901_),
    .Y(_03932_));
 sky130_fd_sc_hd__nand2_1 _08957_ (.A(\core.CPU_Xreg_value_a4[17][28] ),
    .B(_03893_),
    .Y(_03933_));
 sky130_fd_sc_hd__a21oi_1 _08958_ (.A1(_03932_),
    .A2(_03933_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_00868_));
 sky130_fd_sc_hd__nand3_1 _08959_ (.A(\core.CPU_Xreg_value_a4[17][29] ),
    .B(net549),
    .C(net423),
    .Y(_03934_));
 sky130_fd_sc_hd__o21ai_0 _08960_ (.A1(_03523_),
    .A2(net423),
    .B1(_03934_),
    .Y(_00869_));
 sky130_fd_sc_hd__nor2_1 _08961_ (.A(net373),
    .B(net423),
    .Y(_03935_));
 sky130_fd_sc_hd__o21ai_0 _08962_ (.A1(net618),
    .A2(net422),
    .B1(_02644_),
    .Y(_03936_));
 sky130_fd_sc_hd__nor2_1 _08963_ (.A(_03935_),
    .B(_03936_),
    .Y(_00870_));
 sky130_fd_sc_hd__nor2_1 _08964_ (.A(\core.CPU_Xreg_value_a4[17][30] ),
    .B(_03901_),
    .Y(_03937_));
 sky130_fd_sc_hd__a211oi_1 _08965_ (.A1(net345),
    .A2(_03901_),
    .B1(_03937_),
    .C1(net606),
    .Y(_00871_));
 sky130_fd_sc_hd__or3_1 _08966_ (.A(net365),
    .B(net364),
    .C(net423),
    .X(_03938_));
 sky130_fd_sc_hd__nand2_1 _08967_ (.A(\core.CPU_Xreg_value_a4[17][31] ),
    .B(net423),
    .Y(_03939_));
 sky130_fd_sc_hd__a21oi_1 _08968_ (.A1(_03938_),
    .A2(_03939_),
    .B1(net607),
    .Y(_00872_));
 sky130_fd_sc_hd__nand2_1 _08969_ (.A(_03877_),
    .B(net422),
    .Y(_03940_));
 sky130_fd_sc_hd__nand2_1 _08970_ (.A(\core.CPU_Xreg_value_a4[17][3] ),
    .B(net423),
    .Y(_03941_));
 sky130_fd_sc_hd__a21oi_1 _08971_ (.A1(_03940_),
    .A2(_03941_),
    .B1(net607),
    .Y(_00873_));
 sky130_fd_sc_hd__a21oi_1 _08972_ (.A1(net617),
    .A2(net423),
    .B1(net607),
    .Y(_03942_));
 sky130_fd_sc_hd__o21ai_0 _08973_ (.A1(net352),
    .A2(net423),
    .B1(_03942_),
    .Y(_00874_));
 sky130_fd_sc_hd__nand2_1 _08974_ (.A(net371),
    .B(net422),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _08975_ (.A(net616),
    .B(net423),
    .Y(_03944_));
 sky130_fd_sc_hd__a21oi_1 _08976_ (.A1(_03943_),
    .A2(_03944_),
    .B1(net607),
    .Y(_00875_));
 sky130_fd_sc_hd__nand3_1 _08977_ (.A(\core.CPU_Xreg_value_a4[17][6] ),
    .B(_02644_),
    .C(net423),
    .Y(_03945_));
 sky130_fd_sc_hd__o21ai_0 _08978_ (.A1(net344),
    .A2(net423),
    .B1(_03945_),
    .Y(_00876_));
 sky130_fd_sc_hd__o21ai_0 _08979_ (.A1(\core.CPU_Xreg_value_a4[17][7] ),
    .A2(_03901_),
    .B1(net551),
    .Y(_03946_));
 sky130_fd_sc_hd__a21oi_1 _08980_ (.A1(net362),
    .A2(_03901_),
    .B1(_03946_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand3_1 _08981_ (.A(\core.CPU_Xreg_value_a4[17][8] ),
    .B(net551),
    .C(_03893_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_1 _08982_ (.A(net351),
    .B(net422),
    .Y(_03948_));
 sky130_fd_sc_hd__nand2_1 _08983_ (.A(_03947_),
    .B(_03948_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand3_1 _08984_ (.A(\core.CPU_Xreg_value_a4[17][9] ),
    .B(net552),
    .C(_03893_),
    .Y(_03949_));
 sky130_fd_sc_hd__o21ai_0 _08985_ (.A1(_03744_),
    .A2(_03893_),
    .B1(_03949_),
    .Y(_00879_));
 sky130_fd_sc_hd__nor3_1 _08989_ (.A(\core.CPU_rd_a5[3] ),
    .B(\core.CPU_rd_a5[4] ),
    .C(net535),
    .Y(_03953_));
 sky130_fd_sc_hd__a21o_1 _08990_ (.A1(net535),
    .A2(_02554_),
    .B1(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__nand2_2 _08991_ (.A(_03892_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__nand2_1 _08995_ (.A(\core.CPU_Xreg_value_a4[1][0] ),
    .B(_03955_),
    .Y(_03959_));
 sky130_fd_sc_hd__o211ai_1 _08996_ (.A1(_03747_),
    .A2(_03955_),
    .B1(_03959_),
    .C1(net549),
    .Y(_00880_));
 sky130_fd_sc_hd__nand3_1 _08997_ (.A(\core.CPU_Xreg_value_a4[1][10] ),
    .B(net550),
    .C(_03955_),
    .Y(_03960_));
 sky130_fd_sc_hd__o21ai_0 _08998_ (.A1(net348),
    .A2(_03955_),
    .B1(_03960_),
    .Y(_00881_));
 sky130_fd_sc_hd__nand3_1 _08999_ (.A(\core.CPU_Xreg_value_a4[1][11] ),
    .B(net550),
    .C(_03955_),
    .Y(_03961_));
 sky130_fd_sc_hd__o21ai_0 _09000_ (.A1(net361),
    .A2(_03955_),
    .B1(_03961_),
    .Y(_00882_));
 sky130_fd_sc_hd__a21oi_1 _09001_ (.A1(net535),
    .A2(_02554_),
    .B1(_03953_),
    .Y(_03962_));
 sky130_fd_sc_hd__nor2_2 _09002_ (.A(_03900_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__nand2_1 _09004_ (.A(net360),
    .B(net420),
    .Y(_03965_));
 sky130_fd_sc_hd__nand2_1 _09006_ (.A(\core.CPU_Xreg_value_a4[1][12] ),
    .B(net421),
    .Y(_03967_));
 sky130_fd_sc_hd__a21oi_1 _09007_ (.A1(_03965_),
    .A2(_03967_),
    .B1(net606),
    .Y(_00883_));
 sky130_fd_sc_hd__nand3_1 _09008_ (.A(\core.CPU_Xreg_value_a4[1][13] ),
    .B(net552),
    .C(net421),
    .Y(_03968_));
 sky130_fd_sc_hd__o31ai_1 _09009_ (.A1(_02811_),
    .A2(net439),
    .A3(net421),
    .B1(_03968_),
    .Y(_00884_));
 sky130_fd_sc_hd__nand3_1 _09010_ (.A(\core.CPU_Xreg_value_a4[1][14] ),
    .B(net549),
    .C(_03955_),
    .Y(_03969_));
 sky130_fd_sc_hd__o21ai_0 _09011_ (.A1(net347),
    .A2(_03955_),
    .B1(_03969_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand3_1 _09012_ (.A(\core.CPU_Xreg_value_a4[1][15] ),
    .B(net551),
    .C(net421),
    .Y(_03970_));
 sky130_fd_sc_hd__o21ai_0 _09013_ (.A1(_02911_),
    .A2(net421),
    .B1(_03970_),
    .Y(_00886_));
 sky130_fd_sc_hd__o21ai_0 _09016_ (.A1(\core.CPU_Xreg_value_a4[1][16] ),
    .A2(net420),
    .B1(net551),
    .Y(_03973_));
 sky130_fd_sc_hd__a21oi_1 _09017_ (.A1(net346),
    .A2(net420),
    .B1(_03973_),
    .Y(_00887_));
 sky130_fd_sc_hd__nand2_1 _09018_ (.A(_02961_),
    .B(net420),
    .Y(_03974_));
 sky130_fd_sc_hd__nor2_1 _09019_ (.A(_03006_),
    .B(net421),
    .Y(_03975_));
 sky130_fd_sc_hd__a31oi_1 _09020_ (.A1(\core.CPU_Xreg_value_a4[1][17] ),
    .A2(net552),
    .A3(net421),
    .B1(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__o21ai_0 _09021_ (.A1(_03003_),
    .A2(_03974_),
    .B1(_03976_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand3_1 _09022_ (.A(\core.CPU_Xreg_value_a4[1][18] ),
    .B(net552),
    .C(net421),
    .Y(_03977_));
 sky130_fd_sc_hd__o221ai_1 _09023_ (.A1(_03043_),
    .A2(net421),
    .B1(_03974_),
    .B2(net359),
    .C1(_03977_),
    .Y(_00889_));
 sky130_fd_sc_hd__o21ai_0 _09024_ (.A1(\core.CPU_Xreg_value_a4[1][19] ),
    .A2(net420),
    .B1(net551),
    .Y(_03978_));
 sky130_fd_sc_hd__a21oi_1 _09025_ (.A1(net358),
    .A2(net420),
    .B1(_03978_),
    .Y(_00890_));
 sky130_fd_sc_hd__o21ai_0 _09026_ (.A1(\core.CPU_Xreg_value_a4[1][1] ),
    .A2(_03963_),
    .B1(_02644_),
    .Y(_03979_));
 sky130_fd_sc_hd__a21oi_1 _09027_ (.A1(net375),
    .A2(_03963_),
    .B1(_03979_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand3_1 _09028_ (.A(\core.CPU_Xreg_value_a4[1][20] ),
    .B(net549),
    .C(_03955_),
    .Y(_03980_));
 sky130_fd_sc_hd__o21ai_0 _09029_ (.A1(net357),
    .A2(_03955_),
    .B1(_03980_),
    .Y(_00892_));
 sky130_fd_sc_hd__nand3_1 _09030_ (.A(\core.CPU_Xreg_value_a4[1][21] ),
    .B(net550),
    .C(_03955_),
    .Y(_03981_));
 sky130_fd_sc_hd__o21ai_0 _09031_ (.A1(net356),
    .A2(_03955_),
    .B1(_03981_),
    .Y(_00893_));
 sky130_fd_sc_hd__nand2_1 _09032_ (.A(\core.CPU_Xreg_value_a4[1][22] ),
    .B(net421),
    .Y(_03982_));
 sky130_fd_sc_hd__nand2_1 _09033_ (.A(net355),
    .B(net420),
    .Y(_03983_));
 sky130_fd_sc_hd__a21oi_1 _09034_ (.A1(_03982_),
    .A2(_03983_),
    .B1(net607),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2_1 _09035_ (.A(net368),
    .B(net420),
    .Y(_03984_));
 sky130_fd_sc_hd__nand2_1 _09036_ (.A(\core.CPU_Xreg_value_a4[1][23] ),
    .B(net421),
    .Y(_03985_));
 sky130_fd_sc_hd__a21oi_1 _09037_ (.A1(_03984_),
    .A2(_03985_),
    .B1(net606),
    .Y(_00895_));
 sky130_fd_sc_hd__o21ai_0 _09038_ (.A1(\core.CPU_Xreg_value_a4[1][24] ),
    .A2(net420),
    .B1(net551),
    .Y(_03986_));
 sky130_fd_sc_hd__a21oi_2 _09039_ (.A1(_03309_),
    .A2(net420),
    .B1(_03986_),
    .Y(_00896_));
 sky130_fd_sc_hd__o21ai_0 _09040_ (.A1(\core.CPU_Xreg_value_a4[1][25] ),
    .A2(net420),
    .B1(_02644_),
    .Y(_03987_));
 sky130_fd_sc_hd__a21oi_1 _09041_ (.A1(net354),
    .A2(net420),
    .B1(_03987_),
    .Y(_00897_));
 sky130_fd_sc_hd__o21ai_0 _09042_ (.A1(\core.CPU_Xreg_value_a4[1][26] ),
    .A2(net420),
    .B1(net551),
    .Y(_03988_));
 sky130_fd_sc_hd__a21oi_1 _09043_ (.A1(_03389_),
    .A2(net420),
    .B1(_03988_),
    .Y(_00898_));
 sky130_fd_sc_hd__nor2_1 _09044_ (.A(_01114_),
    .B(net421),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2_1 _09045_ (.A(net436),
    .B(net420),
    .Y(_03990_));
 sky130_fd_sc_hd__o21ai_0 _09046_ (.A1(\core.CPU_Xreg_value_a4[1][27] ),
    .A2(net420),
    .B1(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__a311oi_1 _09047_ (.A1(net353),
    .A2(_03431_),
    .A3(_03989_),
    .B1(_03991_),
    .C1(net606),
    .Y(_00899_));
 sky130_fd_sc_hd__nand3_1 _09048_ (.A(_03474_),
    .B(_03475_),
    .C(net420),
    .Y(_03992_));
 sky130_fd_sc_hd__nand2_1 _09049_ (.A(\core.CPU_Xreg_value_a4[1][28] ),
    .B(net421),
    .Y(_03993_));
 sky130_fd_sc_hd__a21oi_1 _09050_ (.A1(_03992_),
    .A2(_03993_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_00900_));
 sky130_fd_sc_hd__nand3_1 _09051_ (.A(\core.CPU_Xreg_value_a4[1][29] ),
    .B(net549),
    .C(_03955_),
    .Y(_03994_));
 sky130_fd_sc_hd__o21ai_0 _09052_ (.A1(_03523_),
    .A2(_03955_),
    .B1(_03994_),
    .Y(_00901_));
 sky130_fd_sc_hd__nor2_1 _09053_ (.A(net373),
    .B(net421),
    .Y(_03995_));
 sky130_fd_sc_hd__o21ai_0 _09054_ (.A1(\core.CPU_Xreg_value_a4[1][2] ),
    .A2(_03963_),
    .B1(_02644_),
    .Y(_03996_));
 sky130_fd_sc_hd__nor2_1 _09055_ (.A(_03995_),
    .B(_03996_),
    .Y(_00902_));
 sky130_fd_sc_hd__o21ai_0 _09056_ (.A1(\core.CPU_Xreg_value_a4[1][30] ),
    .A2(net420),
    .B1(net551),
    .Y(_03997_));
 sky130_fd_sc_hd__a21oi_1 _09057_ (.A1(net345),
    .A2(net420),
    .B1(_03997_),
    .Y(_00903_));
 sky130_fd_sc_hd__or3_1 _09058_ (.A(net365),
    .B(net364),
    .C(_03955_),
    .X(_03998_));
 sky130_fd_sc_hd__nand2_1 _09059_ (.A(\core.CPU_Xreg_value_a4[1][31] ),
    .B(_03955_),
    .Y(_03999_));
 sky130_fd_sc_hd__a21oi_1 _09060_ (.A1(_03998_),
    .A2(_03999_),
    .B1(net607),
    .Y(_00904_));
 sky130_fd_sc_hd__nand2_1 _09061_ (.A(_03877_),
    .B(_03963_),
    .Y(_04000_));
 sky130_fd_sc_hd__nand2_1 _09062_ (.A(\core.CPU_Xreg_value_a4[1][3] ),
    .B(_03955_),
    .Y(_04001_));
 sky130_fd_sc_hd__a21oi_1 _09063_ (.A1(_04000_),
    .A2(_04001_),
    .B1(net607),
    .Y(_00905_));
 sky130_fd_sc_hd__nand3_1 _09065_ (.A(\core.CPU_Xreg_value_a4[1][4] ),
    .B(net549),
    .C(_03955_),
    .Y(_04003_));
 sky130_fd_sc_hd__o21ai_0 _09066_ (.A1(_03662_),
    .A2(_03955_),
    .B1(_04003_),
    .Y(_00906_));
 sky130_fd_sc_hd__nand2_1 _09067_ (.A(net371),
    .B(_03963_),
    .Y(_04004_));
 sky130_fd_sc_hd__nand2_1 _09068_ (.A(\core.CPU_Xreg_value_a4[1][5] ),
    .B(_03955_),
    .Y(_04005_));
 sky130_fd_sc_hd__a21oi_1 _09069_ (.A1(_04004_),
    .A2(_04005_),
    .B1(net607),
    .Y(_00907_));
 sky130_fd_sc_hd__nand3_1 _09070_ (.A(\core.CPU_Xreg_value_a4[1][6] ),
    .B(_02644_),
    .C(net421),
    .Y(_04006_));
 sky130_fd_sc_hd__o21ai_0 _09071_ (.A1(net344),
    .A2(net421),
    .B1(_04006_),
    .Y(_00908_));
 sky130_fd_sc_hd__o21ai_0 _09072_ (.A1(\core.CPU_Xreg_value_a4[1][7] ),
    .A2(net420),
    .B1(net552),
    .Y(_04007_));
 sky130_fd_sc_hd__a21oi_1 _09073_ (.A1(net362),
    .A2(net420),
    .B1(_04007_),
    .Y(_00909_));
 sky130_fd_sc_hd__inv_1 _09074_ (.A(\core.CPU_Xreg_value_a4[1][8] ),
    .Y(_04008_));
 sky130_fd_sc_hd__nand2_1 _09075_ (.A(net351),
    .B(net420),
    .Y(_04009_));
 sky130_fd_sc_hd__o31ai_1 _09076_ (.A1(_04008_),
    .A2(net606),
    .A3(net420),
    .B1(_04009_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand3_1 _09077_ (.A(\core.CPU_Xreg_value_a4[1][9] ),
    .B(net552),
    .C(net421),
    .Y(_04010_));
 sky130_fd_sc_hd__o21ai_0 _09078_ (.A1(_03744_),
    .A2(net421),
    .B1(_04010_),
    .Y(_00911_));
 sky130_fd_sc_hd__and3_1 _09079_ (.A(\core.CPU_rd_a5[3] ),
    .B(\core.CPU_rd_a5[4] ),
    .C(_01114_),
    .X(_04011_));
 sky130_fd_sc_hd__a31oi_1 _09080_ (.A1(\core.CPU_rd_a3[3] ),
    .A2(\core.CPU_rd_a3[4] ),
    .A3(net535),
    .B1(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__a31o_2 _09081_ (.A1(\core.CPU_rd_a3[3] ),
    .A2(\core.CPU_rd_a3[4] ),
    .A3(net535),
    .B1(_04011_),
    .X(_04013_));
 sky130_fd_sc_hd__nor2_2 _09086_ (.A(_02557_),
    .B(_04012_),
    .Y(_04018_));
 sky130_fd_sc_hd__nand2_1 _09088_ (.A(_02545_),
    .B(_04018_),
    .Y(_04020_));
 sky130_fd_sc_hd__nand2_2 _09089_ (.A(_02562_),
    .B(_04013_),
    .Y(_04021_));
 sky130_fd_sc_hd__nand2_1 _09091_ (.A(\core.CPU_Xreg_value_a4[26][0] ),
    .B(net418),
    .Y(_04023_));
 sky130_fd_sc_hd__a21oi_1 _09092_ (.A1(_04020_),
    .A2(_04023_),
    .B1(net607),
    .Y(_00912_));
 sky130_fd_sc_hd__nand3_1 _09095_ (.A(\core.CPU_Xreg_value_a4[26][10] ),
    .B(net550),
    .C(net418),
    .Y(_04026_));
 sky130_fd_sc_hd__o21ai_0 _09096_ (.A1(net348),
    .A2(net418),
    .B1(_04026_),
    .Y(_00913_));
 sky130_fd_sc_hd__nand3_1 _09097_ (.A(\core.CPU_Xreg_value_a4[26][11] ),
    .B(net550),
    .C(net418),
    .Y(_04027_));
 sky130_fd_sc_hd__o21ai_0 _09098_ (.A1(net361),
    .A2(net418),
    .B1(_04027_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_1 _09100_ (.A(\core.CPU_Xreg_value_a4[26][12] ),
    .B(_04021_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _09102_ (.A(net360),
    .B(net419),
    .Y(_04031_));
 sky130_fd_sc_hd__a21oi_1 _09103_ (.A1(_04029_),
    .A2(_04031_),
    .B1(net607),
    .Y(_00915_));
 sky130_fd_sc_hd__nand3_1 _09104_ (.A(\core.CPU_Xreg_value_a4[26][13] ),
    .B(net552),
    .C(_04021_),
    .Y(_04032_));
 sky130_fd_sc_hd__o31ai_1 _09105_ (.A1(_02811_),
    .A2(net439),
    .A3(_04021_),
    .B1(_04032_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand3_1 _09106_ (.A(\core.CPU_Xreg_value_a4[26][14] ),
    .B(net549),
    .C(net418),
    .Y(_04033_));
 sky130_fd_sc_hd__o21ai_0 _09107_ (.A1(net347),
    .A2(net418),
    .B1(_04033_),
    .Y(_00917_));
 sky130_fd_sc_hd__nand3_1 _09108_ (.A(\core.CPU_Xreg_value_a4[26][15] ),
    .B(net551),
    .C(_04021_),
    .Y(_04034_));
 sky130_fd_sc_hd__o21ai_0 _09109_ (.A1(_02911_),
    .A2(_04021_),
    .B1(_04034_),
    .Y(_00918_));
 sky130_fd_sc_hd__o21ai_0 _09110_ (.A1(\core.CPU_Xreg_value_a4[26][16] ),
    .A2(net419),
    .B1(net551),
    .Y(_04035_));
 sky130_fd_sc_hd__a21oi_1 _09111_ (.A1(net346),
    .A2(net419),
    .B1(_04035_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand2_1 _09112_ (.A(_02961_),
    .B(net419),
    .Y(_04036_));
 sky130_fd_sc_hd__nand3_1 _09113_ (.A(\core.CPU_Xreg_value_a4[26][17] ),
    .B(net552),
    .C(_04021_),
    .Y(_04037_));
 sky130_fd_sc_hd__o221ai_1 _09114_ (.A1(_03006_),
    .A2(_04021_),
    .B1(_04036_),
    .B2(_03003_),
    .C1(_04037_),
    .Y(_00920_));
 sky130_fd_sc_hd__nand3_1 _09115_ (.A(\core.CPU_Xreg_value_a4[26][18] ),
    .B(net552),
    .C(_04021_),
    .Y(_04038_));
 sky130_fd_sc_hd__o221ai_1 _09116_ (.A1(_03043_),
    .A2(_04021_),
    .B1(_04036_),
    .B2(net359),
    .C1(_04038_),
    .Y(_00921_));
 sky130_fd_sc_hd__o21ai_0 _09117_ (.A1(\core.CPU_Xreg_value_a4[26][19] ),
    .A2(net419),
    .B1(_02644_),
    .Y(_04039_));
 sky130_fd_sc_hd__a21oi_1 _09118_ (.A1(net358),
    .A2(net419),
    .B1(_04039_),
    .Y(_00922_));
 sky130_fd_sc_hd__nor3_1 _09119_ (.A(\core.CPU_Xreg_value_a4[26][1] ),
    .B(net607),
    .C(_04018_),
    .Y(_04040_));
 sky130_fd_sc_hd__a31oi_1 _09120_ (.A1(_02644_),
    .A2(net375),
    .A3(_04018_),
    .B1(_04040_),
    .Y(_00923_));
 sky130_fd_sc_hd__nand3_1 _09121_ (.A(\core.CPU_Xreg_value_a4[26][20] ),
    .B(net549),
    .C(net418),
    .Y(_04041_));
 sky130_fd_sc_hd__o21ai_0 _09122_ (.A1(net357),
    .A2(net418),
    .B1(_04041_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand3_1 _09123_ (.A(\core.CPU_Xreg_value_a4[26][21] ),
    .B(net550),
    .C(net418),
    .Y(_04042_));
 sky130_fd_sc_hd__o21ai_0 _09124_ (.A1(net356),
    .A2(net418),
    .B1(_04042_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand2_1 _09125_ (.A(\core.CPU_Xreg_value_a4[26][22] ),
    .B(_04021_),
    .Y(_04043_));
 sky130_fd_sc_hd__nand2_1 _09126_ (.A(net355),
    .B(net419),
    .Y(_04044_));
 sky130_fd_sc_hd__a21oi_1 _09127_ (.A1(_04043_),
    .A2(_04044_),
    .B1(net607),
    .Y(_00926_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(net368),
    .B(net419),
    .Y(_04045_));
 sky130_fd_sc_hd__nand2_1 _09129_ (.A(\core.CPU_Xreg_value_a4[26][23] ),
    .B(_04021_),
    .Y(_04046_));
 sky130_fd_sc_hd__a21oi_1 _09130_ (.A1(_04045_),
    .A2(_04046_),
    .B1(net606),
    .Y(_00927_));
 sky130_fd_sc_hd__o21ai_0 _09131_ (.A1(\core.CPU_Xreg_value_a4[26][24] ),
    .A2(net419),
    .B1(net552),
    .Y(_04047_));
 sky130_fd_sc_hd__a21oi_2 _09132_ (.A1(_03309_),
    .A2(net419),
    .B1(_04047_),
    .Y(_00928_));
 sky130_fd_sc_hd__o21ai_0 _09133_ (.A1(\core.CPU_Xreg_value_a4[26][25] ),
    .A2(net419),
    .B1(_02644_),
    .Y(_04048_));
 sky130_fd_sc_hd__a21oi_1 _09134_ (.A1(net354),
    .A2(net419),
    .B1(_04048_),
    .Y(_00929_));
 sky130_fd_sc_hd__o21ai_0 _09135_ (.A1(\core.CPU_Xreg_value_a4[26][26] ),
    .A2(net419),
    .B1(net551),
    .Y(_04049_));
 sky130_fd_sc_hd__a21oi_1 _09136_ (.A1(_03389_),
    .A2(net419),
    .B1(_04049_),
    .Y(_00930_));
 sky130_fd_sc_hd__nor2_1 _09137_ (.A(_01114_),
    .B(_04021_),
    .Y(_04050_));
 sky130_fd_sc_hd__nand2_1 _09138_ (.A(net436),
    .B(net419),
    .Y(_04051_));
 sky130_fd_sc_hd__o21ai_0 _09139_ (.A1(\core.CPU_Xreg_value_a4[26][27] ),
    .A2(net419),
    .B1(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__a311oi_1 _09140_ (.A1(net353),
    .A2(_03431_),
    .A3(_04050_),
    .B1(_04052_),
    .C1(net607),
    .Y(_00931_));
 sky130_fd_sc_hd__nand3_1 _09141_ (.A(_03474_),
    .B(_03475_),
    .C(net419),
    .Y(_04053_));
 sky130_fd_sc_hd__nand2_1 _09142_ (.A(\core.CPU_Xreg_value_a4[26][28] ),
    .B(_04021_),
    .Y(_04054_));
 sky130_fd_sc_hd__a21oi_1 _09143_ (.A1(_04053_),
    .A2(_04054_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_00932_));
 sky130_fd_sc_hd__nand3_1 _09144_ (.A(\core.CPU_Xreg_value_a4[26][29] ),
    .B(net549),
    .C(net418),
    .Y(_04055_));
 sky130_fd_sc_hd__o21ai_0 _09145_ (.A1(_03523_),
    .A2(net418),
    .B1(_04055_),
    .Y(_00933_));
 sky130_fd_sc_hd__nor2_1 _09146_ (.A(net373),
    .B(net418),
    .Y(_04056_));
 sky130_fd_sc_hd__o21ai_0 _09147_ (.A1(\core.CPU_Xreg_value_a4[26][2] ),
    .A2(_04018_),
    .B1(_02644_),
    .Y(_04057_));
 sky130_fd_sc_hd__nor2_1 _09148_ (.A(_04056_),
    .B(_04057_),
    .Y(_00934_));
 sky130_fd_sc_hd__o21ai_0 _09149_ (.A1(\core.CPU_Xreg_value_a4[26][30] ),
    .A2(net419),
    .B1(net551),
    .Y(_04058_));
 sky130_fd_sc_hd__a21oi_1 _09150_ (.A1(net345),
    .A2(net419),
    .B1(_04058_),
    .Y(_00935_));
 sky130_fd_sc_hd__or3_1 _09151_ (.A(net365),
    .B(net364),
    .C(net418),
    .X(_04059_));
 sky130_fd_sc_hd__nand2_1 _09152_ (.A(\core.CPU_Xreg_value_a4[26][31] ),
    .B(net418),
    .Y(_04060_));
 sky130_fd_sc_hd__a21oi_1 _09153_ (.A1(_04059_),
    .A2(_04060_),
    .B1(net607),
    .Y(_00936_));
 sky130_fd_sc_hd__nand2_1 _09154_ (.A(\core.CPU_Xreg_value_a4[26][3] ),
    .B(net418),
    .Y(_04061_));
 sky130_fd_sc_hd__o211ai_1 _09155_ (.A1(net363),
    .A2(net418),
    .B1(_04061_),
    .C1(net549),
    .Y(_00937_));
 sky130_fd_sc_hd__a21oi_1 _09156_ (.A1(\core.CPU_Xreg_value_a4[26][4] ),
    .A2(net418),
    .B1(net607),
    .Y(_04062_));
 sky130_fd_sc_hd__o21ai_0 _09157_ (.A1(net352),
    .A2(net418),
    .B1(_04062_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_1 _09158_ (.A(net371),
    .B(_04018_),
    .Y(_04063_));
 sky130_fd_sc_hd__nand2_1 _09159_ (.A(\core.CPU_Xreg_value_a4[26][5] ),
    .B(net418),
    .Y(_04064_));
 sky130_fd_sc_hd__a21oi_1 _09160_ (.A1(_04063_),
    .A2(_04064_),
    .B1(net607),
    .Y(_00939_));
 sky130_fd_sc_hd__nand3_1 _09161_ (.A(\core.CPU_Xreg_value_a4[26][6] ),
    .B(_02644_),
    .C(net418),
    .Y(_04065_));
 sky130_fd_sc_hd__o21ai_0 _09162_ (.A1(net344),
    .A2(net418),
    .B1(_04065_),
    .Y(_00940_));
 sky130_fd_sc_hd__o21ai_0 _09164_ (.A1(\core.CPU_Xreg_value_a4[26][7] ),
    .A2(net419),
    .B1(net551),
    .Y(_04067_));
 sky130_fd_sc_hd__a21oi_1 _09165_ (.A1(net362),
    .A2(net419),
    .B1(_04067_),
    .Y(_00941_));
 sky130_fd_sc_hd__nand2_1 _09166_ (.A(net351),
    .B(net419),
    .Y(_04068_));
 sky130_fd_sc_hd__nand3_1 _09167_ (.A(\core.CPU_Xreg_value_a4[26][8] ),
    .B(net551),
    .C(_04021_),
    .Y(_04069_));
 sky130_fd_sc_hd__nand2_1 _09168_ (.A(_04068_),
    .B(_04069_),
    .Y(_00942_));
 sky130_fd_sc_hd__nand3_1 _09169_ (.A(\core.CPU_Xreg_value_a4[26][9] ),
    .B(net552),
    .C(_04021_),
    .Y(_04070_));
 sky130_fd_sc_hd__o21ai_0 _09170_ (.A1(_03744_),
    .A2(_04021_),
    .B1(_04070_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand2_2 _09171_ (.A(_03750_),
    .B(_04013_),
    .Y(_04071_));
 sky130_fd_sc_hd__nand2_1 _09175_ (.A(\core.CPU_Xreg_value_a4[27][0] ),
    .B(net417),
    .Y(_04075_));
 sky130_fd_sc_hd__o211ai_1 _09176_ (.A1(_03747_),
    .A2(net417),
    .B1(_04075_),
    .C1(net550),
    .Y(_00944_));
 sky130_fd_sc_hd__nand3_1 _09179_ (.A(\core.CPU_Xreg_value_a4[27][10] ),
    .B(net550),
    .C(net417),
    .Y(_04078_));
 sky130_fd_sc_hd__o21ai_0 _09180_ (.A1(net348),
    .A2(net417),
    .B1(_04078_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand3_1 _09181_ (.A(\core.CPU_Xreg_value_a4[27][11] ),
    .B(net550),
    .C(net417),
    .Y(_04079_));
 sky130_fd_sc_hd__o21ai_0 _09182_ (.A1(net361),
    .A2(net417),
    .B1(_04079_),
    .Y(_00946_));
 sky130_fd_sc_hd__nor2_2 _09183_ (.A(_03760_),
    .B(_04012_),
    .Y(_04080_));
 sky130_fd_sc_hd__nand2_1 _09185_ (.A(net360),
    .B(net416),
    .Y(_04082_));
 sky130_fd_sc_hd__nand2_1 _09186_ (.A(\core.CPU_Xreg_value_a4[27][12] ),
    .B(_04071_),
    .Y(_04083_));
 sky130_fd_sc_hd__a21oi_1 _09188_ (.A1(_04082_),
    .A2(_04083_),
    .B1(net606),
    .Y(_00947_));
 sky130_fd_sc_hd__nand3_1 _09189_ (.A(\core.CPU_Xreg_value_a4[27][13] ),
    .B(net552),
    .C(_04071_),
    .Y(_04085_));
 sky130_fd_sc_hd__o31ai_1 _09190_ (.A1(_02811_),
    .A2(net439),
    .A3(_04071_),
    .B1(_04085_),
    .Y(_00948_));
 sky130_fd_sc_hd__nand3_1 _09191_ (.A(\core.CPU_Xreg_value_a4[27][14] ),
    .B(net549),
    .C(net417),
    .Y(_04086_));
 sky130_fd_sc_hd__o21ai_0 _09192_ (.A1(net347),
    .A2(net417),
    .B1(_04086_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand3_1 _09193_ (.A(\core.CPU_Xreg_value_a4[27][15] ),
    .B(net551),
    .C(net417),
    .Y(_04087_));
 sky130_fd_sc_hd__o21ai_0 _09194_ (.A1(_02911_),
    .A2(net417),
    .B1(_04087_),
    .Y(_00950_));
 sky130_fd_sc_hd__o21ai_0 _09196_ (.A1(\core.CPU_Xreg_value_a4[27][16] ),
    .A2(net416),
    .B1(net551),
    .Y(_04089_));
 sky130_fd_sc_hd__a21oi_1 _09197_ (.A1(net346),
    .A2(net416),
    .B1(_04089_),
    .Y(_00951_));
 sky130_fd_sc_hd__nand2_1 _09198_ (.A(_02961_),
    .B(net416),
    .Y(_04090_));
 sky130_fd_sc_hd__nand3_1 _09199_ (.A(\core.CPU_Xreg_value_a4[27][17] ),
    .B(net552),
    .C(_04071_),
    .Y(_04091_));
 sky130_fd_sc_hd__o221ai_1 _09200_ (.A1(_03006_),
    .A2(_04071_),
    .B1(_04090_),
    .B2(_03003_),
    .C1(_04091_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand3_1 _09201_ (.A(\core.CPU_Xreg_value_a4[27][18] ),
    .B(net552),
    .C(_04071_),
    .Y(_04092_));
 sky130_fd_sc_hd__o221ai_1 _09202_ (.A1(_03043_),
    .A2(_04071_),
    .B1(_04090_),
    .B2(net359),
    .C1(_04092_),
    .Y(_00953_));
 sky130_fd_sc_hd__o21ai_0 _09203_ (.A1(\core.CPU_Xreg_value_a4[27][19] ),
    .A2(net416),
    .B1(_02644_),
    .Y(_04093_));
 sky130_fd_sc_hd__a21oi_1 _09204_ (.A1(net358),
    .A2(net416),
    .B1(_04093_),
    .Y(_00954_));
 sky130_fd_sc_hd__nor3_1 _09205_ (.A(\core.CPU_Xreg_value_a4[27][1] ),
    .B(net607),
    .C(_04080_),
    .Y(_04094_));
 sky130_fd_sc_hd__a31oi_1 _09206_ (.A1(_02644_),
    .A2(net375),
    .A3(_04080_),
    .B1(_04094_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand3_1 _09207_ (.A(\core.CPU_Xreg_value_a4[27][20] ),
    .B(net549),
    .C(net417),
    .Y(_04095_));
 sky130_fd_sc_hd__o21ai_0 _09208_ (.A1(net357),
    .A2(net417),
    .B1(_04095_),
    .Y(_00956_));
 sky130_fd_sc_hd__nand3_1 _09209_ (.A(\core.CPU_Xreg_value_a4[27][21] ),
    .B(net550),
    .C(net417),
    .Y(_04096_));
 sky130_fd_sc_hd__o21ai_0 _09210_ (.A1(net356),
    .A2(net417),
    .B1(_04096_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand2_1 _09211_ (.A(\core.CPU_Xreg_value_a4[27][22] ),
    .B(net417),
    .Y(_04097_));
 sky130_fd_sc_hd__nand2_1 _09212_ (.A(net355),
    .B(net416),
    .Y(_04098_));
 sky130_fd_sc_hd__a21oi_1 _09213_ (.A1(_04097_),
    .A2(_04098_),
    .B1(net607),
    .Y(_00958_));
 sky130_fd_sc_hd__nand2_1 _09214_ (.A(net368),
    .B(net416),
    .Y(_04099_));
 sky130_fd_sc_hd__nand2_1 _09215_ (.A(\core.CPU_Xreg_value_a4[27][23] ),
    .B(net417),
    .Y(_04100_));
 sky130_fd_sc_hd__a21oi_1 _09216_ (.A1(_04099_),
    .A2(_04100_),
    .B1(net606),
    .Y(_00959_));
 sky130_fd_sc_hd__o21ai_0 _09217_ (.A1(\core.CPU_Xreg_value_a4[27][24] ),
    .A2(net416),
    .B1(net552),
    .Y(_04101_));
 sky130_fd_sc_hd__a21oi_2 _09218_ (.A1(_03309_),
    .A2(net416),
    .B1(_04101_),
    .Y(_00960_));
 sky130_fd_sc_hd__o21ai_0 _09219_ (.A1(\core.CPU_Xreg_value_a4[27][25] ),
    .A2(net416),
    .B1(_02644_),
    .Y(_04102_));
 sky130_fd_sc_hd__a21oi_1 _09220_ (.A1(net354),
    .A2(net416),
    .B1(_04102_),
    .Y(_00961_));
 sky130_fd_sc_hd__o21ai_0 _09221_ (.A1(\core.CPU_Xreg_value_a4[27][26] ),
    .A2(net416),
    .B1(net551),
    .Y(_04103_));
 sky130_fd_sc_hd__a21oi_1 _09222_ (.A1(_03389_),
    .A2(net416),
    .B1(_04103_),
    .Y(_00962_));
 sky130_fd_sc_hd__nor2_1 _09223_ (.A(_01114_),
    .B(_04071_),
    .Y(_04104_));
 sky130_fd_sc_hd__nand2_1 _09224_ (.A(net436),
    .B(net416),
    .Y(_04105_));
 sky130_fd_sc_hd__o21ai_0 _09225_ (.A1(\core.CPU_Xreg_value_a4[27][27] ),
    .A2(net416),
    .B1(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__a311oi_1 _09226_ (.A1(net353),
    .A2(_03431_),
    .A3(_04104_),
    .B1(_04106_),
    .C1(net607),
    .Y(_00963_));
 sky130_fd_sc_hd__nand3_1 _09227_ (.A(_03474_),
    .B(_03475_),
    .C(net416),
    .Y(_04107_));
 sky130_fd_sc_hd__nand2_1 _09228_ (.A(\core.CPU_Xreg_value_a4[27][28] ),
    .B(_04071_),
    .Y(_04108_));
 sky130_fd_sc_hd__a21oi_1 _09229_ (.A1(_04107_),
    .A2(_04108_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_00964_));
 sky130_fd_sc_hd__nand3_1 _09230_ (.A(\core.CPU_Xreg_value_a4[27][29] ),
    .B(net549),
    .C(net417),
    .Y(_04109_));
 sky130_fd_sc_hd__o21ai_0 _09231_ (.A1(_03523_),
    .A2(net417),
    .B1(_04109_),
    .Y(_00965_));
 sky130_fd_sc_hd__nor2_1 _09232_ (.A(net373),
    .B(net417),
    .Y(_04110_));
 sky130_fd_sc_hd__o21ai_0 _09233_ (.A1(\core.CPU_Xreg_value_a4[27][2] ),
    .A2(_04080_),
    .B1(_02644_),
    .Y(_04111_));
 sky130_fd_sc_hd__nor2_1 _09234_ (.A(_04110_),
    .B(_04111_),
    .Y(_00966_));
 sky130_fd_sc_hd__o21ai_0 _09235_ (.A1(\core.CPU_Xreg_value_a4[27][30] ),
    .A2(net416),
    .B1(_02644_),
    .Y(_04112_));
 sky130_fd_sc_hd__a21oi_1 _09236_ (.A1(net345),
    .A2(net416),
    .B1(_04112_),
    .Y(_00967_));
 sky130_fd_sc_hd__or3_1 _09237_ (.A(net365),
    .B(net364),
    .C(net417),
    .X(_04113_));
 sky130_fd_sc_hd__nand2_1 _09238_ (.A(\core.CPU_Xreg_value_a4[27][31] ),
    .B(net417),
    .Y(_04114_));
 sky130_fd_sc_hd__a21oi_1 _09239_ (.A1(_04113_),
    .A2(_04114_),
    .B1(net607),
    .Y(_00968_));
 sky130_fd_sc_hd__nand2_1 _09240_ (.A(\core.CPU_Xreg_value_a4[27][3] ),
    .B(net417),
    .Y(_04115_));
 sky130_fd_sc_hd__o211ai_1 _09241_ (.A1(net363),
    .A2(net417),
    .B1(_04115_),
    .C1(net549),
    .Y(_00969_));
 sky130_fd_sc_hd__a21oi_1 _09242_ (.A1(\core.CPU_Xreg_value_a4[27][4] ),
    .A2(net417),
    .B1(net607),
    .Y(_04116_));
 sky130_fd_sc_hd__o21ai_0 _09243_ (.A1(net352),
    .A2(net417),
    .B1(_04116_),
    .Y(_00970_));
 sky130_fd_sc_hd__nand2_1 _09244_ (.A(net371),
    .B(_04080_),
    .Y(_04117_));
 sky130_fd_sc_hd__nand2_1 _09245_ (.A(\core.CPU_Xreg_value_a4[27][5] ),
    .B(net417),
    .Y(_04118_));
 sky130_fd_sc_hd__a21oi_1 _09246_ (.A1(_04117_),
    .A2(_04118_),
    .B1(net607),
    .Y(_00971_));
 sky130_fd_sc_hd__nand3_1 _09247_ (.A(\core.CPU_Xreg_value_a4[27][6] ),
    .B(_02644_),
    .C(net417),
    .Y(_04119_));
 sky130_fd_sc_hd__o21ai_0 _09248_ (.A1(net344),
    .A2(net417),
    .B1(_04119_),
    .Y(_00972_));
 sky130_fd_sc_hd__o21ai_0 _09249_ (.A1(\core.CPU_Xreg_value_a4[27][7] ),
    .A2(net416),
    .B1(net551),
    .Y(_04120_));
 sky130_fd_sc_hd__a21oi_1 _09250_ (.A1(net362),
    .A2(net416),
    .B1(_04120_),
    .Y(_00973_));
 sky130_fd_sc_hd__nand2_1 _09251_ (.A(net351),
    .B(net416),
    .Y(_04121_));
 sky130_fd_sc_hd__nand3_1 _09252_ (.A(\core.CPU_Xreg_value_a4[27][8] ),
    .B(net551),
    .C(net417),
    .Y(_04122_));
 sky130_fd_sc_hd__nand2_1 _09253_ (.A(_04121_),
    .B(_04122_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand3_1 _09254_ (.A(\core.CPU_Xreg_value_a4[27][9] ),
    .B(net552),
    .C(net417),
    .Y(_04123_));
 sky130_fd_sc_hd__o21ai_0 _09255_ (.A1(_03744_),
    .A2(net417),
    .B1(_04123_),
    .Y(_00975_));
 sky130_fd_sc_hd__nor2_4 _09256_ (.A(_02557_),
    .B(_03962_),
    .Y(_04124_));
 sky130_fd_sc_hd__nand2_1 _09258_ (.A(_02545_),
    .B(_04124_),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2_2 _09259_ (.A(_02562_),
    .B(_03954_),
    .Y(_04127_));
 sky130_fd_sc_hd__nand2_1 _09261_ (.A(\core.CPU_Xreg_value_a4[2][0] ),
    .B(_04127_),
    .Y(_04129_));
 sky130_fd_sc_hd__a21oi_1 _09262_ (.A1(_04126_),
    .A2(_04129_),
    .B1(net607),
    .Y(_00976_));
 sky130_fd_sc_hd__nand3_1 _09265_ (.A(\core.CPU_Xreg_value_a4[2][10] ),
    .B(net550),
    .C(_04127_),
    .Y(_04132_));
 sky130_fd_sc_hd__o21ai_0 _09266_ (.A1(net348),
    .A2(_04127_),
    .B1(_04132_),
    .Y(_00977_));
 sky130_fd_sc_hd__nand3_1 _09268_ (.A(\core.CPU_Xreg_value_a4[2][11] ),
    .B(net550),
    .C(_04127_),
    .Y(_04134_));
 sky130_fd_sc_hd__o21ai_0 _09269_ (.A1(net361),
    .A2(_04127_),
    .B1(_04134_),
    .Y(_00978_));
 sky130_fd_sc_hd__nand2_1 _09271_ (.A(net360),
    .B(net415),
    .Y(_04136_));
 sky130_fd_sc_hd__nand2_1 _09272_ (.A(\core.CPU_Xreg_value_a4[2][12] ),
    .B(net414),
    .Y(_04137_));
 sky130_fd_sc_hd__a21oi_1 _09273_ (.A1(_04136_),
    .A2(_04137_),
    .B1(net606),
    .Y(_00979_));
 sky130_fd_sc_hd__nand3_1 _09274_ (.A(\core.CPU_Xreg_value_a4[2][13] ),
    .B(net552),
    .C(net414),
    .Y(_04138_));
 sky130_fd_sc_hd__o31ai_1 _09275_ (.A1(_02811_),
    .A2(net439),
    .A3(net414),
    .B1(_04138_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand3_1 _09276_ (.A(\core.CPU_Xreg_value_a4[2][14] ),
    .B(net549),
    .C(_04127_),
    .Y(_04139_));
 sky130_fd_sc_hd__o21ai_0 _09277_ (.A1(net347),
    .A2(_04127_),
    .B1(_04139_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand3_1 _09278_ (.A(\core.CPU_Xreg_value_a4[2][15] ),
    .B(net551),
    .C(net414),
    .Y(_04140_));
 sky130_fd_sc_hd__o21ai_0 _09279_ (.A1(_02911_),
    .A2(net414),
    .B1(_04140_),
    .Y(_00982_));
 sky130_fd_sc_hd__o21ai_0 _09280_ (.A1(\core.CPU_Xreg_value_a4[2][16] ),
    .A2(net415),
    .B1(net551),
    .Y(_04141_));
 sky130_fd_sc_hd__a21oi_1 _09281_ (.A1(net346),
    .A2(net415),
    .B1(_04141_),
    .Y(_00983_));
 sky130_fd_sc_hd__nand2_1 _09282_ (.A(_02961_),
    .B(net415),
    .Y(_04142_));
 sky130_fd_sc_hd__nand3_1 _09283_ (.A(\core.CPU_Xreg_value_a4[2][17] ),
    .B(net552),
    .C(net414),
    .Y(_04143_));
 sky130_fd_sc_hd__o221ai_1 _09284_ (.A1(_03006_),
    .A2(net414),
    .B1(_04142_),
    .B2(_03003_),
    .C1(_04143_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand3_1 _09285_ (.A(\core.CPU_Xreg_value_a4[2][18] ),
    .B(net552),
    .C(net414),
    .Y(_04144_));
 sky130_fd_sc_hd__o221ai_1 _09286_ (.A1(_03043_),
    .A2(net414),
    .B1(_04142_),
    .B2(net359),
    .C1(_04144_),
    .Y(_00985_));
 sky130_fd_sc_hd__o21ai_0 _09287_ (.A1(\core.CPU_Xreg_value_a4[2][19] ),
    .A2(net415),
    .B1(_02644_),
    .Y(_04145_));
 sky130_fd_sc_hd__a21oi_1 _09288_ (.A1(net358),
    .A2(net415),
    .B1(_04145_),
    .Y(_00986_));
 sky130_fd_sc_hd__nor2_1 _09289_ (.A(net607),
    .B(net414),
    .Y(_04146_));
 sky130_fd_sc_hd__nor3_1 _09290_ (.A(\core.CPU_Xreg_value_a4[2][1] ),
    .B(net607),
    .C(_04124_),
    .Y(_04147_));
 sky130_fd_sc_hd__a21oi_1 _09291_ (.A1(net375),
    .A2(_04146_),
    .B1(_04147_),
    .Y(_00987_));
 sky130_fd_sc_hd__nand3_1 _09292_ (.A(\core.CPU_Xreg_value_a4[2][20] ),
    .B(net549),
    .C(_04127_),
    .Y(_04148_));
 sky130_fd_sc_hd__o21ai_0 _09293_ (.A1(net357),
    .A2(_04127_),
    .B1(_04148_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand3_1 _09294_ (.A(\core.CPU_Xreg_value_a4[2][21] ),
    .B(net550),
    .C(_04127_),
    .Y(_04149_));
 sky130_fd_sc_hd__o21ai_0 _09295_ (.A1(net356),
    .A2(_04127_),
    .B1(_04149_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_1 _09296_ (.A(\core.CPU_Xreg_value_a4[2][22] ),
    .B(net414),
    .Y(_04150_));
 sky130_fd_sc_hd__nand2_1 _09297_ (.A(net355),
    .B(net415),
    .Y(_04151_));
 sky130_fd_sc_hd__a21oi_1 _09298_ (.A1(_04150_),
    .A2(_04151_),
    .B1(net607),
    .Y(_00990_));
 sky130_fd_sc_hd__nand2_1 _09299_ (.A(net368),
    .B(net415),
    .Y(_04152_));
 sky130_fd_sc_hd__nand2_1 _09300_ (.A(\core.CPU_Xreg_value_a4[2][23] ),
    .B(net414),
    .Y(_04153_));
 sky130_fd_sc_hd__a21oi_1 _09301_ (.A1(_04152_),
    .A2(_04153_),
    .B1(net606),
    .Y(_00991_));
 sky130_fd_sc_hd__o21ai_0 _09303_ (.A1(\core.CPU_Xreg_value_a4[2][24] ),
    .A2(net415),
    .B1(net551),
    .Y(_04155_));
 sky130_fd_sc_hd__a21oi_1 _09304_ (.A1(_03309_),
    .A2(net415),
    .B1(_04155_),
    .Y(_00992_));
 sky130_fd_sc_hd__o21ai_0 _09305_ (.A1(\core.CPU_Xreg_value_a4[2][25] ),
    .A2(net415),
    .B1(_02644_),
    .Y(_04156_));
 sky130_fd_sc_hd__a21oi_1 _09306_ (.A1(net354),
    .A2(net415),
    .B1(_04156_),
    .Y(_00993_));
 sky130_fd_sc_hd__o21ai_0 _09307_ (.A1(\core.CPU_Xreg_value_a4[2][26] ),
    .A2(net415),
    .B1(net551),
    .Y(_04157_));
 sky130_fd_sc_hd__a21oi_1 _09308_ (.A1(_03389_),
    .A2(net415),
    .B1(_04157_),
    .Y(_00994_));
 sky130_fd_sc_hd__nor2_1 _09309_ (.A(_01114_),
    .B(net414),
    .Y(_04158_));
 sky130_fd_sc_hd__nand2_1 _09310_ (.A(net436),
    .B(net415),
    .Y(_04159_));
 sky130_fd_sc_hd__o21ai_0 _09311_ (.A1(\core.CPU_Xreg_value_a4[2][27] ),
    .A2(net415),
    .B1(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__a311oi_1 _09312_ (.A1(net353),
    .A2(_03431_),
    .A3(_04158_),
    .B1(_04160_),
    .C1(net606),
    .Y(_00995_));
 sky130_fd_sc_hd__nand3_1 _09313_ (.A(_03474_),
    .B(_03475_),
    .C(net415),
    .Y(_04161_));
 sky130_fd_sc_hd__nand2_1 _09314_ (.A(\core.CPU_Xreg_value_a4[2][28] ),
    .B(net414),
    .Y(_04162_));
 sky130_fd_sc_hd__a21oi_1 _09316_ (.A1(_04161_),
    .A2(_04162_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_00996_));
 sky130_fd_sc_hd__inv_1 _09317_ (.A(\core.CPU_Xreg_value_a4[2][29] ),
    .Y(_04164_));
 sky130_fd_sc_hd__nand2_1 _09318_ (.A(net366),
    .B(_04146_),
    .Y(_04165_));
 sky130_fd_sc_hd__o31ai_1 _09319_ (.A1(_04164_),
    .A2(net607),
    .A3(_04124_),
    .B1(_04165_),
    .Y(_00997_));
 sky130_fd_sc_hd__nor2_1 _09320_ (.A(net373),
    .B(net414),
    .Y(_04166_));
 sky130_fd_sc_hd__o21ai_0 _09321_ (.A1(\core.CPU_Xreg_value_a4[2][2] ),
    .A2(_04124_),
    .B1(_02644_),
    .Y(_04167_));
 sky130_fd_sc_hd__nor2_1 _09322_ (.A(_04166_),
    .B(_04167_),
    .Y(_00998_));
 sky130_fd_sc_hd__o21ai_0 _09323_ (.A1(\core.CPU_Xreg_value_a4[2][30] ),
    .A2(net415),
    .B1(net551),
    .Y(_04168_));
 sky130_fd_sc_hd__a21oi_1 _09324_ (.A1(net345),
    .A2(net415),
    .B1(_04168_),
    .Y(_00999_));
 sky130_fd_sc_hd__or3_1 _09325_ (.A(net365),
    .B(net364),
    .C(_04127_),
    .X(_04169_));
 sky130_fd_sc_hd__nand2_1 _09326_ (.A(\core.CPU_Xreg_value_a4[2][31] ),
    .B(net414),
    .Y(_04170_));
 sky130_fd_sc_hd__a21oi_1 _09327_ (.A1(_04169_),
    .A2(_04170_),
    .B1(net607),
    .Y(_01000_));
 sky130_fd_sc_hd__nand2_1 _09328_ (.A(_03877_),
    .B(_04124_),
    .Y(_04171_));
 sky130_fd_sc_hd__nand2_1 _09329_ (.A(\core.CPU_Xreg_value_a4[2][3] ),
    .B(_04127_),
    .Y(_04172_));
 sky130_fd_sc_hd__a21oi_1 _09330_ (.A1(_04171_),
    .A2(_04172_),
    .B1(net607),
    .Y(_01001_));
 sky130_fd_sc_hd__nand3_1 _09331_ (.A(\core.CPU_Xreg_value_a4[2][4] ),
    .B(net549),
    .C(_04127_),
    .Y(_04173_));
 sky130_fd_sc_hd__o21ai_0 _09332_ (.A1(_03662_),
    .A2(_04127_),
    .B1(_04173_),
    .Y(_01002_));
 sky130_fd_sc_hd__nand2_1 _09333_ (.A(net371),
    .B(_04124_),
    .Y(_04174_));
 sky130_fd_sc_hd__nand2_1 _09334_ (.A(\core.CPU_Xreg_value_a4[2][5] ),
    .B(_04127_),
    .Y(_04175_));
 sky130_fd_sc_hd__a21oi_1 _09335_ (.A1(_04174_),
    .A2(_04175_),
    .B1(net607),
    .Y(_01003_));
 sky130_fd_sc_hd__nand3_1 _09336_ (.A(\core.CPU_Xreg_value_a4[2][6] ),
    .B(_02644_),
    .C(net414),
    .Y(_04176_));
 sky130_fd_sc_hd__o21ai_0 _09337_ (.A1(net344),
    .A2(net414),
    .B1(_04176_),
    .Y(_01004_));
 sky130_fd_sc_hd__o21ai_0 _09338_ (.A1(\core.CPU_Xreg_value_a4[2][7] ),
    .A2(net415),
    .B1(net552),
    .Y(_04177_));
 sky130_fd_sc_hd__a21oi_1 _09339_ (.A1(net362),
    .A2(net415),
    .B1(_04177_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_1 _09340_ (.A(net351),
    .B(net415),
    .Y(_04178_));
 sky130_fd_sc_hd__nand3_1 _09341_ (.A(\core.CPU_Xreg_value_a4[2][8] ),
    .B(net551),
    .C(net414),
    .Y(_04179_));
 sky130_fd_sc_hd__nand2_1 _09342_ (.A(_04178_),
    .B(_04179_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand3_1 _09343_ (.A(\core.CPU_Xreg_value_a4[2][9] ),
    .B(net552),
    .C(net414),
    .Y(_04180_));
 sky130_fd_sc_hd__o21ai_0 _09344_ (.A1(_03744_),
    .A2(net414),
    .B1(_04180_),
    .Y(_01007_));
 sky130_fd_sc_hd__nand2_2 _09345_ (.A(_03750_),
    .B(_03954_),
    .Y(_04181_));
 sky130_fd_sc_hd__nand2_1 _09349_ (.A(\core.CPU_Xreg_value_a4[3][0] ),
    .B(net413),
    .Y(_04185_));
 sky130_fd_sc_hd__o211ai_1 _09350_ (.A1(_03747_),
    .A2(net413),
    .B1(_04185_),
    .C1(net549),
    .Y(_01008_));
 sky130_fd_sc_hd__nand3_1 _09351_ (.A(\core.CPU_Xreg_value_a4[3][10] ),
    .B(net550),
    .C(net413),
    .Y(_04186_));
 sky130_fd_sc_hd__o21ai_0 _09352_ (.A1(net348),
    .A2(net413),
    .B1(_04186_),
    .Y(_01009_));
 sky130_fd_sc_hd__nand3_1 _09353_ (.A(\core.CPU_Xreg_value_a4[3][11] ),
    .B(net550),
    .C(net413),
    .Y(_04187_));
 sky130_fd_sc_hd__o21ai_0 _09354_ (.A1(net361),
    .A2(net413),
    .B1(_04187_),
    .Y(_01010_));
 sky130_fd_sc_hd__nor2_2 _09355_ (.A(_03760_),
    .B(_03962_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand2_1 _09357_ (.A(net360),
    .B(net412),
    .Y(_04190_));
 sky130_fd_sc_hd__nand2_1 _09359_ (.A(\core.CPU_Xreg_value_a4[3][12] ),
    .B(_04181_),
    .Y(_04192_));
 sky130_fd_sc_hd__a21oi_1 _09360_ (.A1(_04190_),
    .A2(_04192_),
    .B1(net607),
    .Y(_01011_));
 sky130_fd_sc_hd__nand3_1 _09361_ (.A(\core.CPU_Xreg_value_a4[3][13] ),
    .B(net552),
    .C(_04181_),
    .Y(_04193_));
 sky130_fd_sc_hd__o31ai_1 _09362_ (.A1(_02811_),
    .A2(net439),
    .A3(_04181_),
    .B1(_04193_),
    .Y(_01012_));
 sky130_fd_sc_hd__nand3_1 _09364_ (.A(\core.CPU_Xreg_value_a4[3][14] ),
    .B(net549),
    .C(net413),
    .Y(_04195_));
 sky130_fd_sc_hd__o21ai_0 _09365_ (.A1(net347),
    .A2(net413),
    .B1(_04195_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand3_1 _09366_ (.A(\core.CPU_Xreg_value_a4[3][15] ),
    .B(net551),
    .C(_04181_),
    .Y(_04196_));
 sky130_fd_sc_hd__o21ai_0 _09367_ (.A1(_02911_),
    .A2(_04181_),
    .B1(_04196_),
    .Y(_01014_));
 sky130_fd_sc_hd__o21ai_0 _09369_ (.A1(\core.CPU_Xreg_value_a4[3][16] ),
    .A2(net412),
    .B1(net551),
    .Y(_04198_));
 sky130_fd_sc_hd__a21oi_1 _09370_ (.A1(net346),
    .A2(net412),
    .B1(_04198_),
    .Y(_01015_));
 sky130_fd_sc_hd__nand2_1 _09371_ (.A(_02961_),
    .B(net412),
    .Y(_04199_));
 sky130_fd_sc_hd__nor2_1 _09372_ (.A(_03006_),
    .B(_04181_),
    .Y(_04200_));
 sky130_fd_sc_hd__a31oi_1 _09373_ (.A1(\core.CPU_Xreg_value_a4[3][17] ),
    .A2(net551),
    .A3(_04181_),
    .B1(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__o21ai_0 _09374_ (.A1(_03003_),
    .A2(_04199_),
    .B1(_04201_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand3_1 _09375_ (.A(\core.CPU_Xreg_value_a4[3][18] ),
    .B(net552),
    .C(_04181_),
    .Y(_04202_));
 sky130_fd_sc_hd__o221ai_1 _09376_ (.A1(_03043_),
    .A2(_04181_),
    .B1(_04199_),
    .B2(net359),
    .C1(_04202_),
    .Y(_01017_));
 sky130_fd_sc_hd__o21ai_0 _09377_ (.A1(\core.CPU_Xreg_value_a4[3][19] ),
    .A2(net412),
    .B1(_02644_),
    .Y(_04203_));
 sky130_fd_sc_hd__a21oi_1 _09378_ (.A1(net358),
    .A2(net412),
    .B1(_04203_),
    .Y(_01018_));
 sky130_fd_sc_hd__nor3_1 _09379_ (.A(\core.CPU_Xreg_value_a4[3][1] ),
    .B(net607),
    .C(_04188_),
    .Y(_04204_));
 sky130_fd_sc_hd__a31oi_1 _09380_ (.A1(net549),
    .A2(net375),
    .A3(_04188_),
    .B1(_04204_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand3_1 _09381_ (.A(\core.CPU_Xreg_value_a4[3][20] ),
    .B(net549),
    .C(net413),
    .Y(_04205_));
 sky130_fd_sc_hd__o21ai_0 _09382_ (.A1(net357),
    .A2(net413),
    .B1(_04205_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand3_1 _09383_ (.A(\core.CPU_Xreg_value_a4[3][21] ),
    .B(net550),
    .C(net413),
    .Y(_04206_));
 sky130_fd_sc_hd__o21ai_0 _09384_ (.A1(net356),
    .A2(net413),
    .B1(_04206_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _09385_ (.A(\core.CPU_Xreg_value_a4[3][22] ),
    .B(_04181_),
    .Y(_04207_));
 sky130_fd_sc_hd__nand2_1 _09386_ (.A(net355),
    .B(net412),
    .Y(_04208_));
 sky130_fd_sc_hd__a21oi_1 _09387_ (.A1(_04207_),
    .A2(_04208_),
    .B1(net606),
    .Y(_01022_));
 sky130_fd_sc_hd__nand2_1 _09388_ (.A(net368),
    .B(net412),
    .Y(_04209_));
 sky130_fd_sc_hd__nand2_1 _09389_ (.A(\core.CPU_Xreg_value_a4[3][23] ),
    .B(_04181_),
    .Y(_04210_));
 sky130_fd_sc_hd__a21oi_1 _09390_ (.A1(_04209_),
    .A2(_04210_),
    .B1(net606),
    .Y(_01023_));
 sky130_fd_sc_hd__o21ai_0 _09391_ (.A1(\core.CPU_Xreg_value_a4[3][24] ),
    .A2(net412),
    .B1(net552),
    .Y(_04211_));
 sky130_fd_sc_hd__a21oi_1 _09392_ (.A1(_03309_),
    .A2(net412),
    .B1(_04211_),
    .Y(_01024_));
 sky130_fd_sc_hd__o21ai_0 _09393_ (.A1(\core.CPU_Xreg_value_a4[3][25] ),
    .A2(net412),
    .B1(_02644_),
    .Y(_04212_));
 sky130_fd_sc_hd__a21oi_1 _09394_ (.A1(net354),
    .A2(net412),
    .B1(_04212_),
    .Y(_01025_));
 sky130_fd_sc_hd__o21ai_0 _09395_ (.A1(\core.CPU_Xreg_value_a4[3][26] ),
    .A2(net412),
    .B1(net551),
    .Y(_04213_));
 sky130_fd_sc_hd__a21oi_1 _09396_ (.A1(_03389_),
    .A2(net412),
    .B1(_04213_),
    .Y(_01026_));
 sky130_fd_sc_hd__nor2_1 _09397_ (.A(_01114_),
    .B(_04181_),
    .Y(_04214_));
 sky130_fd_sc_hd__nand2_1 _09398_ (.A(net436),
    .B(net412),
    .Y(_04215_));
 sky130_fd_sc_hd__o21ai_0 _09399_ (.A1(\core.CPU_Xreg_value_a4[3][27] ),
    .A2(net412),
    .B1(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__a311oi_1 _09400_ (.A1(net353),
    .A2(_03431_),
    .A3(_04214_),
    .B1(_04216_),
    .C1(net606),
    .Y(_01027_));
 sky130_fd_sc_hd__nand3_1 _09401_ (.A(_03474_),
    .B(_03475_),
    .C(net412),
    .Y(_04217_));
 sky130_fd_sc_hd__nand2_1 _09402_ (.A(\core.CPU_Xreg_value_a4[3][28] ),
    .B(_04181_),
    .Y(_04218_));
 sky130_fd_sc_hd__a21oi_1 _09403_ (.A1(_04217_),
    .A2(_04218_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_01028_));
 sky130_fd_sc_hd__nand3_1 _09404_ (.A(\core.CPU_Xreg_value_a4[3][29] ),
    .B(net549),
    .C(net413),
    .Y(_04219_));
 sky130_fd_sc_hd__o21ai_0 _09405_ (.A1(_03523_),
    .A2(net413),
    .B1(_04219_),
    .Y(_01029_));
 sky130_fd_sc_hd__nor2_1 _09406_ (.A(net373),
    .B(net413),
    .Y(_04220_));
 sky130_fd_sc_hd__o21ai_0 _09407_ (.A1(\core.CPU_Xreg_value_a4[3][2] ),
    .A2(_04188_),
    .B1(_02644_),
    .Y(_04221_));
 sky130_fd_sc_hd__nor2_1 _09408_ (.A(_04220_),
    .B(_04221_),
    .Y(_01030_));
 sky130_fd_sc_hd__o21ai_0 _09410_ (.A1(\core.CPU_Xreg_value_a4[3][30] ),
    .A2(net412),
    .B1(net551),
    .Y(_04223_));
 sky130_fd_sc_hd__a21oi_1 _09411_ (.A1(net345),
    .A2(net412),
    .B1(_04223_),
    .Y(_01031_));
 sky130_fd_sc_hd__or3_1 _09412_ (.A(net365),
    .B(net364),
    .C(net413),
    .X(_04224_));
 sky130_fd_sc_hd__nand2_1 _09413_ (.A(\core.CPU_Xreg_value_a4[3][31] ),
    .B(net413),
    .Y(_04225_));
 sky130_fd_sc_hd__a21oi_1 _09414_ (.A1(_04224_),
    .A2(_04225_),
    .B1(net607),
    .Y(_01032_));
 sky130_fd_sc_hd__nand2_1 _09415_ (.A(_03877_),
    .B(_04188_),
    .Y(_04226_));
 sky130_fd_sc_hd__nand2_1 _09416_ (.A(\core.CPU_Xreg_value_a4[3][3] ),
    .B(net413),
    .Y(_04227_));
 sky130_fd_sc_hd__a21oi_1 _09417_ (.A1(_04226_),
    .A2(_04227_),
    .B1(net607),
    .Y(_01033_));
 sky130_fd_sc_hd__nand3_1 _09418_ (.A(\core.CPU_Xreg_value_a4[3][4] ),
    .B(net549),
    .C(net413),
    .Y(_04228_));
 sky130_fd_sc_hd__o21ai_0 _09419_ (.A1(_03662_),
    .A2(net413),
    .B1(_04228_),
    .Y(_01034_));
 sky130_fd_sc_hd__nand2_1 _09420_ (.A(net371),
    .B(_04188_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand2_1 _09421_ (.A(\core.CPU_Xreg_value_a4[3][5] ),
    .B(net413),
    .Y(_04230_));
 sky130_fd_sc_hd__a21oi_1 _09423_ (.A1(_04229_),
    .A2(_04230_),
    .B1(net607),
    .Y(_01035_));
 sky130_fd_sc_hd__nand3_1 _09424_ (.A(\core.CPU_Xreg_value_a4[3][6] ),
    .B(_02644_),
    .C(net413),
    .Y(_04232_));
 sky130_fd_sc_hd__o21ai_0 _09425_ (.A1(net344),
    .A2(net413),
    .B1(_04232_),
    .Y(_01036_));
 sky130_fd_sc_hd__o21ai_0 _09426_ (.A1(\core.CPU_Xreg_value_a4[3][7] ),
    .A2(net412),
    .B1(net552),
    .Y(_04233_));
 sky130_fd_sc_hd__a21oi_1 _09427_ (.A1(net362),
    .A2(net412),
    .B1(_04233_),
    .Y(_01037_));
 sky130_fd_sc_hd__nand2_1 _09428_ (.A(net351),
    .B(net412),
    .Y(_04234_));
 sky130_fd_sc_hd__nand3_1 _09429_ (.A(\core.CPU_Xreg_value_a4[3][8] ),
    .B(net551),
    .C(_04181_),
    .Y(_04235_));
 sky130_fd_sc_hd__nand2_1 _09430_ (.A(_04234_),
    .B(_04235_),
    .Y(_01038_));
 sky130_fd_sc_hd__nand3_1 _09431_ (.A(\core.CPU_Xreg_value_a4[3][9] ),
    .B(net552),
    .C(_04181_),
    .Y(_04236_));
 sky130_fd_sc_hd__o21ai_0 _09432_ (.A1(_03744_),
    .A2(_04181_),
    .B1(_04236_),
    .Y(_01039_));
 sky130_fd_sc_hd__nor3_2 _09433_ (.A(_02550_),
    .B(_03825_),
    .C(_03830_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_1 _09435_ (.A(_02545_),
    .B(net411),
    .Y(_04239_));
 sky130_fd_sc_hd__nand2_2 _09436_ (.A(_02561_),
    .B(_03835_),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2_1 _09438_ (.A(\core.CPU_Xreg_value_a4[8][0] ),
    .B(net389),
    .Y(_04242_));
 sky130_fd_sc_hd__a21oi_1 _09439_ (.A1(_04239_),
    .A2(_04242_),
    .B1(net607),
    .Y(_01040_));
 sky130_fd_sc_hd__nand3_1 _09442_ (.A(\core.CPU_Xreg_value_a4[8][10] ),
    .B(net550),
    .C(net389),
    .Y(_04245_));
 sky130_fd_sc_hd__o21ai_0 _09443_ (.A1(net348),
    .A2(net389),
    .B1(_04245_),
    .Y(_01041_));
 sky130_fd_sc_hd__nand3_1 _09444_ (.A(\core.CPU_Xreg_value_a4[8][11] ),
    .B(net550),
    .C(net389),
    .Y(_04246_));
 sky130_fd_sc_hd__o21ai_0 _09445_ (.A1(net361),
    .A2(net389),
    .B1(_04246_),
    .Y(_01042_));
 sky130_fd_sc_hd__nand2_1 _09447_ (.A(net360),
    .B(net411),
    .Y(_04248_));
 sky130_fd_sc_hd__nand2_1 _09448_ (.A(\core.CPU_Xreg_value_a4[8][12] ),
    .B(net389),
    .Y(_04249_));
 sky130_fd_sc_hd__a21oi_1 _09449_ (.A1(_04248_),
    .A2(_04249_),
    .B1(net607),
    .Y(_01043_));
 sky130_fd_sc_hd__nand3_1 _09450_ (.A(\core.CPU_Xreg_value_a4[8][13] ),
    .B(net552),
    .C(net389),
    .Y(_04250_));
 sky130_fd_sc_hd__o31ai_1 _09451_ (.A1(_02811_),
    .A2(net439),
    .A3(net389),
    .B1(_04250_),
    .Y(_01044_));
 sky130_fd_sc_hd__nand3_1 _09454_ (.A(\core.CPU_Xreg_value_a4[8][14] ),
    .B(net549),
    .C(net389),
    .Y(_04253_));
 sky130_fd_sc_hd__o21ai_0 _09455_ (.A1(net347),
    .A2(net389),
    .B1(_04253_),
    .Y(_01045_));
 sky130_fd_sc_hd__nand3_1 _09456_ (.A(\core.CPU_Xreg_value_a4[8][15] ),
    .B(net551),
    .C(net389),
    .Y(_04254_));
 sky130_fd_sc_hd__o21ai_0 _09457_ (.A1(_02911_),
    .A2(net389),
    .B1(_04254_),
    .Y(_01046_));
 sky130_fd_sc_hd__o21ai_0 _09458_ (.A1(\core.CPU_Xreg_value_a4[8][16] ),
    .A2(net411),
    .B1(net551),
    .Y(_04255_));
 sky130_fd_sc_hd__a21oi_1 _09459_ (.A1(net346),
    .A2(net411),
    .B1(_04255_),
    .Y(_01047_));
 sky130_fd_sc_hd__nand2_1 _09460_ (.A(_02961_),
    .B(net411),
    .Y(_04256_));
 sky130_fd_sc_hd__nand3_1 _09461_ (.A(\core.CPU_Xreg_value_a4[8][17] ),
    .B(net551),
    .C(net389),
    .Y(_04257_));
 sky130_fd_sc_hd__o221ai_1 _09462_ (.A1(_03006_),
    .A2(net389),
    .B1(_04256_),
    .B2(_03003_),
    .C1(_04257_),
    .Y(_01048_));
 sky130_fd_sc_hd__nand3_1 _09463_ (.A(\core.CPU_Xreg_value_a4[8][18] ),
    .B(net552),
    .C(net389),
    .Y(_04258_));
 sky130_fd_sc_hd__o221ai_1 _09464_ (.A1(_03043_),
    .A2(net389),
    .B1(_04256_),
    .B2(net359),
    .C1(_04258_),
    .Y(_01049_));
 sky130_fd_sc_hd__o21ai_0 _09465_ (.A1(\core.CPU_Xreg_value_a4[8][19] ),
    .A2(net411),
    .B1(net551),
    .Y(_04259_));
 sky130_fd_sc_hd__a21oi_1 _09466_ (.A1(net358),
    .A2(net411),
    .B1(_04259_),
    .Y(_01050_));
 sky130_fd_sc_hd__o21ai_0 _09467_ (.A1(\core.CPU_Xreg_value_a4[8][1] ),
    .A2(net411),
    .B1(_02644_),
    .Y(_04260_));
 sky130_fd_sc_hd__a21oi_1 _09468_ (.A1(net375),
    .A2(net411),
    .B1(_04260_),
    .Y(_01051_));
 sky130_fd_sc_hd__nand3_1 _09469_ (.A(\core.CPU_Xreg_value_a4[8][20] ),
    .B(net550),
    .C(net389),
    .Y(_04261_));
 sky130_fd_sc_hd__o21ai_0 _09470_ (.A1(net357),
    .A2(net389),
    .B1(_04261_),
    .Y(_01052_));
 sky130_fd_sc_hd__nand3_1 _09471_ (.A(\core.CPU_Xreg_value_a4[8][21] ),
    .B(net550),
    .C(net389),
    .Y(_04262_));
 sky130_fd_sc_hd__o21ai_0 _09472_ (.A1(net356),
    .A2(net389),
    .B1(_04262_),
    .Y(_01053_));
 sky130_fd_sc_hd__nand2_1 _09473_ (.A(\core.CPU_Xreg_value_a4[8][22] ),
    .B(net389),
    .Y(_04263_));
 sky130_fd_sc_hd__nand2_1 _09474_ (.A(net355),
    .B(net411),
    .Y(_04264_));
 sky130_fd_sc_hd__a21oi_1 _09475_ (.A1(_04263_),
    .A2(_04264_),
    .B1(net607),
    .Y(_01054_));
 sky130_fd_sc_hd__nand2_1 _09476_ (.A(net368),
    .B(net411),
    .Y(_04265_));
 sky130_fd_sc_hd__nand2_1 _09477_ (.A(\core.CPU_Xreg_value_a4[8][23] ),
    .B(net389),
    .Y(_04266_));
 sky130_fd_sc_hd__a21oi_1 _09478_ (.A1(_04265_),
    .A2(_04266_),
    .B1(net606),
    .Y(_01055_));
 sky130_fd_sc_hd__o21ai_0 _09479_ (.A1(\core.CPU_Xreg_value_a4[8][24] ),
    .A2(net411),
    .B1(net552),
    .Y(_04267_));
 sky130_fd_sc_hd__a21oi_1 _09480_ (.A1(_03309_),
    .A2(net411),
    .B1(_04267_),
    .Y(_01056_));
 sky130_fd_sc_hd__o21ai_0 _09481_ (.A1(\core.CPU_Xreg_value_a4[8][25] ),
    .A2(net411),
    .B1(_02644_),
    .Y(_04268_));
 sky130_fd_sc_hd__a21oi_1 _09482_ (.A1(net354),
    .A2(net411),
    .B1(_04268_),
    .Y(_01057_));
 sky130_fd_sc_hd__o21ai_0 _09483_ (.A1(\core.CPU_Xreg_value_a4[8][26] ),
    .A2(net411),
    .B1(net551),
    .Y(_04269_));
 sky130_fd_sc_hd__a21oi_1 _09484_ (.A1(_03389_),
    .A2(net411),
    .B1(_04269_),
    .Y(_01058_));
 sky130_fd_sc_hd__nor2_1 _09485_ (.A(_01114_),
    .B(net389),
    .Y(_04270_));
 sky130_fd_sc_hd__nand2_1 _09486_ (.A(net436),
    .B(net411),
    .Y(_04271_));
 sky130_fd_sc_hd__o21ai_0 _09487_ (.A1(\core.CPU_Xreg_value_a4[8][27] ),
    .A2(net411),
    .B1(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__a311oi_1 _09488_ (.A1(net353),
    .A2(_03431_),
    .A3(_04270_),
    .B1(_04272_),
    .C1(net606),
    .Y(_01059_));
 sky130_fd_sc_hd__nand3_1 _09489_ (.A(_03474_),
    .B(_03475_),
    .C(net411),
    .Y(_04273_));
 sky130_fd_sc_hd__nand2_1 _09490_ (.A(\core.CPU_Xreg_value_a4[8][28] ),
    .B(net389),
    .Y(_04274_));
 sky130_fd_sc_hd__a21oi_1 _09491_ (.A1(_04273_),
    .A2(_04274_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_01060_));
 sky130_fd_sc_hd__nand3_1 _09492_ (.A(\core.CPU_Xreg_value_a4[8][29] ),
    .B(net549),
    .C(net389),
    .Y(_04275_));
 sky130_fd_sc_hd__o21ai_0 _09493_ (.A1(_03523_),
    .A2(net389),
    .B1(_04275_),
    .Y(_01061_));
 sky130_fd_sc_hd__nor2_1 _09494_ (.A(net373),
    .B(net389),
    .Y(_04276_));
 sky130_fd_sc_hd__o21ai_0 _09495_ (.A1(\core.CPU_Xreg_value_a4[8][2] ),
    .A2(net411),
    .B1(_02644_),
    .Y(_04277_));
 sky130_fd_sc_hd__nor2_1 _09496_ (.A(_04276_),
    .B(_04277_),
    .Y(_01062_));
 sky130_fd_sc_hd__o21ai_0 _09497_ (.A1(\core.CPU_Xreg_value_a4[8][30] ),
    .A2(net411),
    .B1(_02644_),
    .Y(_04278_));
 sky130_fd_sc_hd__a21oi_1 _09498_ (.A1(net345),
    .A2(net411),
    .B1(_04278_),
    .Y(_01063_));
 sky130_fd_sc_hd__or3_1 _09499_ (.A(net365),
    .B(net364),
    .C(net389),
    .X(_04279_));
 sky130_fd_sc_hd__nand2_1 _09500_ (.A(\core.CPU_Xreg_value_a4[8][31] ),
    .B(net389),
    .Y(_04280_));
 sky130_fd_sc_hd__a21oi_1 _09501_ (.A1(_04279_),
    .A2(_04280_),
    .B1(net607),
    .Y(_01064_));
 sky130_fd_sc_hd__nand2_1 _09502_ (.A(\core.CPU_Xreg_value_a4[8][3] ),
    .B(net389),
    .Y(_04281_));
 sky130_fd_sc_hd__o211ai_1 _09503_ (.A1(net363),
    .A2(net389),
    .B1(_04281_),
    .C1(net549),
    .Y(_01065_));
 sky130_fd_sc_hd__nand3_1 _09504_ (.A(\core.CPU_Xreg_value_a4[8][4] ),
    .B(net549),
    .C(net389),
    .Y(_04282_));
 sky130_fd_sc_hd__o21ai_0 _09505_ (.A1(_03662_),
    .A2(net389),
    .B1(_04282_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand2_1 _09506_ (.A(net371),
    .B(net411),
    .Y(_04283_));
 sky130_fd_sc_hd__nand2_1 _09507_ (.A(\core.CPU_Xreg_value_a4[8][5] ),
    .B(net389),
    .Y(_04284_));
 sky130_fd_sc_hd__a21oi_1 _09508_ (.A1(_04283_),
    .A2(_04284_),
    .B1(net607),
    .Y(_01067_));
 sky130_fd_sc_hd__nand3_1 _09509_ (.A(\core.CPU_Xreg_value_a4[8][6] ),
    .B(_02644_),
    .C(net389),
    .Y(_04285_));
 sky130_fd_sc_hd__o21ai_0 _09510_ (.A1(net344),
    .A2(net389),
    .B1(_04285_),
    .Y(_01068_));
 sky130_fd_sc_hd__o21ai_0 _09511_ (.A1(\core.CPU_Xreg_value_a4[8][7] ),
    .A2(net411),
    .B1(net552),
    .Y(_04286_));
 sky130_fd_sc_hd__a21oi_1 _09512_ (.A1(net362),
    .A2(net411),
    .B1(_04286_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand2_1 _09513_ (.A(net351),
    .B(net411),
    .Y(_04287_));
 sky130_fd_sc_hd__nand3_1 _09514_ (.A(\core.CPU_Xreg_value_a4[8][8] ),
    .B(net551),
    .C(net389),
    .Y(_04288_));
 sky130_fd_sc_hd__nand2_1 _09515_ (.A(_04287_),
    .B(_04288_),
    .Y(_01070_));
 sky130_fd_sc_hd__nand3_1 _09516_ (.A(\core.CPU_Xreg_value_a4[8][9] ),
    .B(net552),
    .C(net389),
    .Y(_04289_));
 sky130_fd_sc_hd__o21ai_0 _09517_ (.A1(_03744_),
    .A2(net389),
    .B1(_04289_),
    .Y(_01071_));
 sky130_fd_sc_hd__nand2_2 _09518_ (.A(_02561_),
    .B(_03892_),
    .Y(_04290_));
 sky130_fd_sc_hd__nand2_1 _09522_ (.A(\core.CPU_Xreg_value_a4[9][0] ),
    .B(net410),
    .Y(_04294_));
 sky130_fd_sc_hd__o211ai_1 _09523_ (.A1(_03747_),
    .A2(net410),
    .B1(_04294_),
    .C1(net549),
    .Y(_01072_));
 sky130_fd_sc_hd__nand3_1 _09524_ (.A(\core.CPU_Xreg_value_a4[9][10] ),
    .B(net550),
    .C(net410),
    .Y(_04295_));
 sky130_fd_sc_hd__o21ai_0 _09525_ (.A1(net348),
    .A2(net410),
    .B1(_04295_),
    .Y(_01073_));
 sky130_fd_sc_hd__nand3_1 _09527_ (.A(\core.CPU_Xreg_value_a4[9][11] ),
    .B(net550),
    .C(net410),
    .Y(_04297_));
 sky130_fd_sc_hd__o21ai_0 _09528_ (.A1(net361),
    .A2(net410),
    .B1(_04297_),
    .Y(_01074_));
 sky130_fd_sc_hd__nor2_2 _09529_ (.A(_02550_),
    .B(_03900_),
    .Y(_04298_));
 sky130_fd_sc_hd__nand2_1 _09531_ (.A(net360),
    .B(net409),
    .Y(_04300_));
 sky130_fd_sc_hd__nand2_1 _09532_ (.A(\core.CPU_Xreg_value_a4[9][12] ),
    .B(_04290_),
    .Y(_04301_));
 sky130_fd_sc_hd__a21oi_1 _09533_ (.A1(_04300_),
    .A2(_04301_),
    .B1(net607),
    .Y(_01075_));
 sky130_fd_sc_hd__nand3_1 _09534_ (.A(\core.CPU_Xreg_value_a4[9][13] ),
    .B(net552),
    .C(_04290_),
    .Y(_04302_));
 sky130_fd_sc_hd__o31ai_1 _09535_ (.A1(_02811_),
    .A2(net439),
    .A3(_04290_),
    .B1(_04302_),
    .Y(_01076_));
 sky130_fd_sc_hd__nand3_1 _09536_ (.A(\core.CPU_Xreg_value_a4[9][14] ),
    .B(net549),
    .C(net410),
    .Y(_04303_));
 sky130_fd_sc_hd__o21ai_0 _09537_ (.A1(net347),
    .A2(net410),
    .B1(_04303_),
    .Y(_01077_));
 sky130_fd_sc_hd__nand3_1 _09538_ (.A(\core.CPU_Xreg_value_a4[9][15] ),
    .B(net551),
    .C(_04290_),
    .Y(_04304_));
 sky130_fd_sc_hd__o21ai_0 _09539_ (.A1(_02911_),
    .A2(_04290_),
    .B1(_04304_),
    .Y(_01078_));
 sky130_fd_sc_hd__o21ai_0 _09541_ (.A1(\core.CPU_Xreg_value_a4[9][16] ),
    .A2(net409),
    .B1(net551),
    .Y(_04306_));
 sky130_fd_sc_hd__a21oi_1 _09542_ (.A1(net346),
    .A2(net409),
    .B1(_04306_),
    .Y(_01079_));
 sky130_fd_sc_hd__nand2_1 _09543_ (.A(_02961_),
    .B(net409),
    .Y(_04307_));
 sky130_fd_sc_hd__nor2_1 _09544_ (.A(_03006_),
    .B(_04290_),
    .Y(_04308_));
 sky130_fd_sc_hd__a31oi_1 _09545_ (.A1(\core.CPU_Xreg_value_a4[9][17] ),
    .A2(net551),
    .A3(_04290_),
    .B1(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__o21ai_0 _09546_ (.A1(_03003_),
    .A2(_04307_),
    .B1(_04309_),
    .Y(_01080_));
 sky130_fd_sc_hd__nand3_1 _09547_ (.A(\core.CPU_Xreg_value_a4[9][18] ),
    .B(net552),
    .C(_04290_),
    .Y(_04310_));
 sky130_fd_sc_hd__o221ai_1 _09548_ (.A1(_03043_),
    .A2(_04290_),
    .B1(_04307_),
    .B2(net359),
    .C1(_04310_),
    .Y(_01081_));
 sky130_fd_sc_hd__o21ai_0 _09549_ (.A1(\core.CPU_Xreg_value_a4[9][19] ),
    .A2(net409),
    .B1(_02644_),
    .Y(_04311_));
 sky130_fd_sc_hd__a21oi_1 _09550_ (.A1(net358),
    .A2(net409),
    .B1(_04311_),
    .Y(_01082_));
 sky130_fd_sc_hd__o21ai_0 _09551_ (.A1(\core.CPU_Xreg_value_a4[9][1] ),
    .A2(net409),
    .B1(_02644_),
    .Y(_04312_));
 sky130_fd_sc_hd__a21oi_1 _09552_ (.A1(net375),
    .A2(net409),
    .B1(_04312_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand3_1 _09553_ (.A(\core.CPU_Xreg_value_a4[9][20] ),
    .B(net550),
    .C(net410),
    .Y(_04313_));
 sky130_fd_sc_hd__o21ai_0 _09554_ (.A1(net357),
    .A2(net410),
    .B1(_04313_),
    .Y(_01084_));
 sky130_fd_sc_hd__nand3_1 _09555_ (.A(\core.CPU_Xreg_value_a4[9][21] ),
    .B(net550),
    .C(net410),
    .Y(_04314_));
 sky130_fd_sc_hd__o21ai_0 _09556_ (.A1(net356),
    .A2(net410),
    .B1(_04314_),
    .Y(_01085_));
 sky130_fd_sc_hd__nand2_1 _09557_ (.A(\core.CPU_Xreg_value_a4[9][22] ),
    .B(_04290_),
    .Y(_04315_));
 sky130_fd_sc_hd__nand2_1 _09558_ (.A(net355),
    .B(net409),
    .Y(_04316_));
 sky130_fd_sc_hd__a21oi_1 _09559_ (.A1(_04315_),
    .A2(_04316_),
    .B1(net606),
    .Y(_01086_));
 sky130_fd_sc_hd__nand2_1 _09560_ (.A(net368),
    .B(net409),
    .Y(_04317_));
 sky130_fd_sc_hd__nand2_1 _09561_ (.A(\core.CPU_Xreg_value_a4[9][23] ),
    .B(_04290_),
    .Y(_04318_));
 sky130_fd_sc_hd__a21oi_1 _09562_ (.A1(_04317_),
    .A2(_04318_),
    .B1(net606),
    .Y(_01087_));
 sky130_fd_sc_hd__o21ai_0 _09563_ (.A1(\core.CPU_Xreg_value_a4[9][24] ),
    .A2(net409),
    .B1(net552),
    .Y(_04319_));
 sky130_fd_sc_hd__a21oi_1 _09564_ (.A1(_03309_),
    .A2(net409),
    .B1(_04319_),
    .Y(_01088_));
 sky130_fd_sc_hd__o21ai_0 _09565_ (.A1(\core.CPU_Xreg_value_a4[9][25] ),
    .A2(net409),
    .B1(_02644_),
    .Y(_04320_));
 sky130_fd_sc_hd__a21oi_1 _09566_ (.A1(net354),
    .A2(net409),
    .B1(_04320_),
    .Y(_01089_));
 sky130_fd_sc_hd__o21ai_0 _09567_ (.A1(\core.CPU_Xreg_value_a4[9][26] ),
    .A2(net409),
    .B1(net551),
    .Y(_04321_));
 sky130_fd_sc_hd__a21oi_1 _09568_ (.A1(_03389_),
    .A2(net409),
    .B1(_04321_),
    .Y(_01090_));
 sky130_fd_sc_hd__nor2_1 _09569_ (.A(_01114_),
    .B(_04290_),
    .Y(_04322_));
 sky130_fd_sc_hd__nand2_1 _09570_ (.A(net436),
    .B(net409),
    .Y(_04323_));
 sky130_fd_sc_hd__o21ai_0 _09571_ (.A1(\core.CPU_Xreg_value_a4[9][27] ),
    .A2(net409),
    .B1(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__a311oi_1 _09572_ (.A1(net353),
    .A2(_03431_),
    .A3(_04322_),
    .B1(_04324_),
    .C1(net606),
    .Y(_01091_));
 sky130_fd_sc_hd__nand3_1 _09573_ (.A(_03474_),
    .B(_03475_),
    .C(net409),
    .Y(_04325_));
 sky130_fd_sc_hd__nand2_1 _09574_ (.A(\core.CPU_Xreg_value_a4[9][28] ),
    .B(_04290_),
    .Y(_04326_));
 sky130_fd_sc_hd__a21oi_1 _09575_ (.A1(_04325_),
    .A2(_04326_),
    .B1(\core.CPU_reset_a3 ),
    .Y(_01092_));
 sky130_fd_sc_hd__nand3_1 _09576_ (.A(\core.CPU_Xreg_value_a4[9][29] ),
    .B(net549),
    .C(net410),
    .Y(_04327_));
 sky130_fd_sc_hd__o21ai_0 _09577_ (.A1(_03523_),
    .A2(net410),
    .B1(_04327_),
    .Y(_01093_));
 sky130_fd_sc_hd__nor2_1 _09578_ (.A(net373),
    .B(net410),
    .Y(_04328_));
 sky130_fd_sc_hd__o21ai_0 _09579_ (.A1(\core.CPU_Xreg_value_a4[9][2] ),
    .A2(net409),
    .B1(_02644_),
    .Y(_04329_));
 sky130_fd_sc_hd__nor2_1 _09580_ (.A(_04328_),
    .B(_04329_),
    .Y(_01094_));
 sky130_fd_sc_hd__o21ai_0 _09581_ (.A1(\core.CPU_Xreg_value_a4[9][30] ),
    .A2(net409),
    .B1(_02644_),
    .Y(_04330_));
 sky130_fd_sc_hd__a21oi_1 _09582_ (.A1(net345),
    .A2(net409),
    .B1(_04330_),
    .Y(_01095_));
 sky130_fd_sc_hd__or3_1 _09583_ (.A(net365),
    .B(net364),
    .C(net410),
    .X(_04331_));
 sky130_fd_sc_hd__nand2_1 _09584_ (.A(\core.CPU_Xreg_value_a4[9][31] ),
    .B(net410),
    .Y(_04332_));
 sky130_fd_sc_hd__a21oi_1 _09585_ (.A1(_04331_),
    .A2(_04332_),
    .B1(net607),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(\core.CPU_Xreg_value_a4[9][3] ),
    .B(net410),
    .Y(_04333_));
 sky130_fd_sc_hd__o211ai_1 _09587_ (.A1(net363),
    .A2(net410),
    .B1(_04333_),
    .C1(net549),
    .Y(_01097_));
 sky130_fd_sc_hd__nand3_1 _09588_ (.A(\core.CPU_Xreg_value_a4[9][4] ),
    .B(net549),
    .C(net410),
    .Y(_04334_));
 sky130_fd_sc_hd__o21ai_0 _09589_ (.A1(_03662_),
    .A2(net410),
    .B1(_04334_),
    .Y(_01098_));
 sky130_fd_sc_hd__nand2_1 _09590_ (.A(net371),
    .B(net409),
    .Y(_04335_));
 sky130_fd_sc_hd__nand2_1 _09591_ (.A(\core.CPU_Xreg_value_a4[9][5] ),
    .B(net410),
    .Y(_04336_));
 sky130_fd_sc_hd__a21oi_1 _09592_ (.A1(_04335_),
    .A2(_04336_),
    .B1(net607),
    .Y(_01099_));
 sky130_fd_sc_hd__nand3_1 _09593_ (.A(\core.CPU_Xreg_value_a4[9][6] ),
    .B(_02644_),
    .C(net410),
    .Y(_04337_));
 sky130_fd_sc_hd__o21ai_0 _09594_ (.A1(net344),
    .A2(net410),
    .B1(_04337_),
    .Y(_01100_));
 sky130_fd_sc_hd__o21ai_0 _09595_ (.A1(\core.CPU_Xreg_value_a4[9][7] ),
    .A2(net409),
    .B1(net552),
    .Y(_04338_));
 sky130_fd_sc_hd__a21oi_1 _09596_ (.A1(net362),
    .A2(net409),
    .B1(_04338_),
    .Y(_01101_));
 sky130_fd_sc_hd__nand2_1 _09597_ (.A(net351),
    .B(net409),
    .Y(_04339_));
 sky130_fd_sc_hd__nand3_1 _09598_ (.A(\core.CPU_Xreg_value_a4[9][8] ),
    .B(net551),
    .C(_04290_),
    .Y(_04340_));
 sky130_fd_sc_hd__nand2_1 _09599_ (.A(_04339_),
    .B(_04340_),
    .Y(_01102_));
 sky130_fd_sc_hd__nand3_1 _09600_ (.A(\core.CPU_Xreg_value_a4[9][9] ),
    .B(net552),
    .C(_04290_),
    .Y(_04341_));
 sky130_fd_sc_hd__o21ai_0 _09601_ (.A1(_03744_),
    .A2(_04290_),
    .B1(_04341_),
    .Y(_01103_));
 sky130_fd_sc_hd__nand2_1 _09602_ (.A(\core.CPU_br_tgt_pc_a3[2] ),
    .B(net377),
    .Y(_04342_));
 sky130_fd_sc_hd__nand2_1 _09603_ (.A(\core.CPU_imem_rd_addr_a1[0] ),
    .B(_01168_),
    .Y(_04343_));
 sky130_fd_sc_hd__o221ai_1 _09604_ (.A1(net562),
    .A2(_01166_),
    .B1(_01168_),
    .B2(\core.CPU_inc_pc_a3[2] ),
    .C1(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__a21oi_1 _09605_ (.A1(_04342_),
    .A2(_04344_),
    .B1(net608),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _09606_ (.A(\core.CPU_inc_pc_a3[3] ),
    .B(\core.CPU_valid_load_a3 ),
    .Y(_04345_));
 sky130_fd_sc_hd__nand2_1 _09607_ (.A(\core.CPU_inc_pc_a1[3] ),
    .B(_01168_),
    .Y(_04346_));
 sky130_fd_sc_hd__a21oi_1 _09608_ (.A1(_04345_),
    .A2(_04346_),
    .B1(net377),
    .Y(_04347_));
 sky130_fd_sc_hd__a21oi_1 _09609_ (.A1(\core.CPU_br_tgt_pc_a3[3] ),
    .A2(net377),
    .B1(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__nor2_1 _09610_ (.A(net608),
    .B(_04348_),
    .Y(_01105_));
 sky130_fd_sc_hd__mux2i_1 _09611_ (.A0(\core.CPU_inc_pc_a3[4] ),
    .A1(\core.CPU_inc_pc_a1[4] ),
    .S(_01168_),
    .Y(_04349_));
 sky130_fd_sc_hd__nand2_1 _09612_ (.A(\core.CPU_br_tgt_pc_a3[4] ),
    .B(net377),
    .Y(_04350_));
 sky130_fd_sc_hd__o21ai_0 _09613_ (.A1(net377),
    .A2(_04349_),
    .B1(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__nor2b_1 _09614_ (.A(net608),
    .B_N(_04351_),
    .Y(_01106_));
 sky130_fd_sc_hd__mux2i_1 _09615_ (.A0(\core.CPU_inc_pc_a3[5] ),
    .A1(\core.CPU_inc_pc_a1[5] ),
    .S(_01168_),
    .Y(_04352_));
 sky130_fd_sc_hd__nand2_1 _09616_ (.A(\core.CPU_br_tgt_pc_a3[5] ),
    .B(net377),
    .Y(_04353_));
 sky130_fd_sc_hd__o21ai_0 _09617_ (.A1(net377),
    .A2(_04352_),
    .B1(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__nor2b_1 _09618_ (.A(net608),
    .B_N(_04354_),
    .Y(_01107_));
 sky130_fd_sc_hd__nor2_1 _09619_ (.A(_00204_),
    .B(_00207_),
    .Y(_04355_));
 sky130_fd_sc_hd__nand3b_1 _09620_ (.A_N(_00206_),
    .B(_04355_),
    .C(_00205_),
    .Y(_04356_));
 sky130_fd_sc_hd__nand2b_1 _09621_ (.A_N(net615),
    .B(net614),
    .Y(_04357_));
 sky130_fd_sc_hd__nand2_1 _09622_ (.A(\core.CPU_imem_rd_addr_a1[3] ),
    .B(_00204_),
    .Y(_04358_));
 sky130_fd_sc_hd__o21ai_0 _09623_ (.A1(\core.CPU_imem_rd_addr_a1[3] ),
    .A2(_04356_),
    .B1(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__nand2_1 _09624_ (.A(net615),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__o21ai_0 _09625_ (.A1(_04356_),
    .A2(_04357_),
    .B1(_04360_),
    .Y(\core.CPU_imm_a1[10] ));
 sky130_fd_sc_hd__and2_1 _09626_ (.A(\core.CPU_imem_rd_data_a1[11] ),
    .B(\core.CPU_imm_a1[10] ),
    .X(_01108_));
 sky130_fd_sc_hd__nand2_1 _09627_ (.A(\core.CPU_inc_pc_a3[0] ),
    .B(\core.CPU_valid_load_a3 ),
    .Y(_04361_));
 sky130_fd_sc_hd__nand2_1 _09628_ (.A(\core.CPU_inc_pc_a1[0] ),
    .B(_01168_),
    .Y(_04362_));
 sky130_fd_sc_hd__a21oi_1 _09629_ (.A1(_04361_),
    .A2(_04362_),
    .B1(net377),
    .Y(_04363_));
 sky130_fd_sc_hd__a21oi_1 _09630_ (.A1(\core.CPU_br_tgt_pc_a3[0] ),
    .A2(net377),
    .B1(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__nor2_1 _09631_ (.A(net608),
    .B(_04364_),
    .Y(_01109_));
 sky130_fd_sc_hd__nand2_1 _09632_ (.A(\core.CPU_inc_pc_a3[1] ),
    .B(\core.CPU_valid_load_a3 ),
    .Y(_04365_));
 sky130_fd_sc_hd__nand2_1 _09633_ (.A(\core.CPU_inc_pc_a1[1] ),
    .B(_01168_),
    .Y(_04366_));
 sky130_fd_sc_hd__a21oi_1 _09634_ (.A1(_04365_),
    .A2(_04366_),
    .B1(net377),
    .Y(_04367_));
 sky130_fd_sc_hd__a21oi_1 _09635_ (.A1(\core.CPU_br_tgt_pc_a3[1] ),
    .A2(net377),
    .B1(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__nor2_1 _09636_ (.A(net608),
    .B(_04368_),
    .Y(_01110_));
 sky130_fd_sc_hd__xnor2_1 _09637_ (.A(net615),
    .B(\core.CPU_imem_rd_addr_a1[3] ),
    .Y(_04369_));
 sky130_fd_sc_hd__a21oi_1 _09638_ (.A1(_01183_),
    .A2(_04355_),
    .B1(_04369_),
    .Y(_01111_));
 sky130_fd_sc_hd__nor2_1 _09639_ (.A(_01183_),
    .B(_04369_),
    .Y(_01112_));
 sky130_fd_sc_hd__nor2_1 _09640_ (.A(_04355_),
    .B(_04369_),
    .Y(_01113_));
 sky130_fd_sc_hd__xnor2_1 _09641_ (.A(\core.CPU_pc_a2[2] ),
    .B(_00013_),
    .Y(\core.CPU_br_tgt_pc_a2[2] ));
 sky130_fd_sc_hd__a21o_1 _09642_ (.A1(_00202_),
    .A2(_00016_),
    .B1(_00015_),
    .X(_04370_));
 sky130_fd_sc_hd__nand2_1 _09643_ (.A(\core.CPU_pc_a2[2] ),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__xnor2_1 _09644_ (.A(_00018_),
    .B(_04371_),
    .Y(\core.CPU_br_tgt_pc_a2[3] ));
 sky130_fd_sc_hd__inv_1 _09645_ (.A(_00013_),
    .Y(_04372_));
 sky130_fd_sc_hd__a31oi_1 _09646_ (.A1(\core.CPU_pc_a2[2] ),
    .A2(_04372_),
    .A3(_00018_),
    .B1(_00017_),
    .Y(_04373_));
 sky130_fd_sc_hd__xnor2_1 _09647_ (.A(_00020_),
    .B(_04373_),
    .Y(\core.CPU_br_tgt_pc_a2[4] ));
 sky130_fd_sc_hd__a31o_2 _09648_ (.A1(\core.CPU_pc_a2[2] ),
    .A2(_00018_),
    .A3(_04370_),
    .B1(_00017_),
    .X(_04374_));
 sky130_fd_sc_hd__a21oi_1 _09649_ (.A1(_00020_),
    .A2(_04374_),
    .B1(_00019_),
    .Y(_04375_));
 sky130_fd_sc_hd__xor2_1 _09650_ (.A(\core.CPU_pc_a2[5] ),
    .B(\core.CPU_imm_a2[5] ),
    .X(_04376_));
 sky130_fd_sc_hd__xnor2_1 _09651_ (.A(_04375_),
    .B(_04376_),
    .Y(\core.CPU_br_tgt_pc_a2[5] ));
 sky130_fd_sc_hd__nor2_1 _09652_ (.A(_00205_),
    .B(_00207_),
    .Y(_04377_));
 sky130_fd_sc_hd__nor3_1 _09653_ (.A(net614),
    .B(_00206_),
    .C(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__nand3b_1 _09654_ (.A_N(\core.CPU_imem_rd_addr_a1[3] ),
    .B(_04356_),
    .C(net615),
    .Y(_04379_));
 sky130_fd_sc_hd__o21ai_0 _09655_ (.A1(net615),
    .A2(_04378_),
    .B1(_04379_),
    .Y(\core.CPU_imem_rd_data_a1[20] ));
 sky130_fd_sc_hd__o21a_1 _09656_ (.A1(_00206_),
    .A2(_00204_),
    .B1(net614),
    .X(_04380_));
 sky130_fd_sc_hd__o22ai_1 _09657_ (.A1(net614),
    .A2(_00204_),
    .B1(_04380_),
    .B2(net615),
    .Y(_04381_));
 sky130_fd_sc_hd__nor2_1 _09658_ (.A(net615),
    .B(_01179_),
    .Y(\core.CPU_imm_a1[1] ));
 sky130_fd_sc_hd__a21o_1 _09659_ (.A1(_04377_),
    .A2(_04381_),
    .B1(\core.CPU_imm_a1[1] ),
    .X(\core.CPU_imm_a1[0] ));
 sky130_fd_sc_hd__o21ai_0 _09660_ (.A1(_04356_),
    .A2(_04357_),
    .B1(_04360_),
    .Y(\core.CPU_imm_a1[11] ));
 sky130_fd_sc_hd__mux2i_1 _09661_ (.A0(_00206_),
    .A1(_00205_),
    .S(net615),
    .Y(_04382_));
 sky130_fd_sc_hd__o22ai_1 _09662_ (.A1(_04355_),
    .A2(_04369_),
    .B1(_04382_),
    .B2(\core.CPU_imem_rd_addr_a1[3] ),
    .Y(\core.CPU_imem_rd_data_a1[21] ));
 sky130_fd_sc_hd__o21ai_0 _09663_ (.A1(_04356_),
    .A2(_04357_),
    .B1(_04360_),
    .Y(\core.CPU_imm_a1[12] ));
 sky130_fd_sc_hd__a211oi_1 _09664_ (.A1(\core.CPU_imem_rd_addr_a1[3] ),
    .A2(_00205_),
    .B1(_00206_),
    .C1(net615),
    .Y(_04383_));
 sky130_fd_sc_hd__a21oi_1 _09665_ (.A1(net615),
    .A2(_01181_),
    .B1(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__or2_2 _09666_ (.A(_01113_),
    .B(_04384_),
    .X(\core.CPU_imem_rd_data_a1[23] ));
 sky130_fd_sc_hd__or2_2 _09667_ (.A(_01108_),
    .B(\core.CPU_imm_a1[1] ),
    .X(\core.CPU_imm_a1[3] ));
 sky130_fd_sc_hd__nor3_1 _09668_ (.A(_00206_),
    .B(_00204_),
    .C(_00207_),
    .Y(_04385_));
 sky130_fd_sc_hd__nand3_1 _09669_ (.A(net614),
    .B(_00205_),
    .C(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__nand2_1 _09670_ (.A(_01179_),
    .B(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__mux2_2 _09671_ (.A0(_04387_),
    .A1(_04359_),
    .S(net615),
    .X(\core.CPU_imm_a1[5] ));
 sky130_fd_sc_hd__nor4b_1 _09672_ (.A(\core.CPU_imem_rd_addr_a1[3] ),
    .B(_00205_),
    .C(_04355_),
    .D_N(net615),
    .Y(\core.CPU_is_add_a1 ));
 sky130_fd_sc_hd__o41a_1 _09673_ (.A1(_00205_),
    .A2(_00206_),
    .A3(_00204_),
    .A4(_00207_),
    .B1(net614),
    .X(_04388_));
 sky130_fd_sc_hd__nor2_1 _09674_ (.A(net614),
    .B(_00204_),
    .Y(_04389_));
 sky130_fd_sc_hd__nand2_1 _09675_ (.A(_04377_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__o21ai_0 _09676_ (.A1(net615),
    .A2(_04388_),
    .B1(_04390_),
    .Y(\core.CPU_is_addi_a1 ));
 sky130_fd_sc_hd__and3_1 _09677_ (.A(\core.CPU_imem_rd_addr_a1[2] ),
    .B(net614),
    .C(_00204_),
    .X(\core.CPU_is_beq_a1 ));
 sky130_fd_sc_hd__and2_1 _09678_ (.A(\core.CPU_imem_rd_data_a1[11] ),
    .B(\core.CPU_imm_a1[10] ),
    .X(\core.CPU_is_bne_a1 ));
 sky130_fd_sc_hd__nor3_1 _09679_ (.A(_00205_),
    .B(_04385_),
    .C(_04357_),
    .Y(\core.CPU_is_sub_a1 ));
 sky130_fd_sc_hd__a21oi_1 _09680_ (.A1(\core.CPU_imem_rd_addr_a1[3] ),
    .A2(_00205_),
    .B1(net615),
    .Y(_04391_));
 sky130_fd_sc_hd__a31o_2 _09681_ (.A1(net615),
    .A2(_01181_),
    .A3(_04358_),
    .B1(_04391_),
    .X(\core.CPU_rd_valid_a1 ));
 sky130_fd_sc_hd__inv_1 _09682_ (.A(_03535_),
    .Y(\core.CPU_result_a3[2] ));
 sky130_fd_sc_hd__inv_1 _09683_ (.A(_03659_),
    .Y(\core.CPU_result_a3[4] ));
 sky130_fd_sc_hd__inv_1 _09684_ (.A(_03675_),
    .Y(\core.CPU_result_a3[5] ));
 sky130_fd_sc_hd__nand3_1 _09686_ (.A(\core.CPU_rd_a3[1] ),
    .B(\core.CPU_rd_a3[3] ),
    .C(net595),
    .Y(_04393_));
 sky130_fd_sc_hd__or3_1 _09687_ (.A(\core.CPU_rd_a3[1] ),
    .B(\core.CPU_rd_a3[3] ),
    .C(net595),
    .X(_04394_));
 sky130_fd_sc_hd__xor2_1 _09689_ (.A(\core.CPU_rd_a3[0] ),
    .B(\core.CPU_rf_rd_index1_a2[0] ),
    .X(_04396_));
 sky130_fd_sc_hd__xor2_1 _09691_ (.A(\core.CPU_rd_a3[4] ),
    .B(\core.CPU_rf_rd_index1_a2[4] ),
    .X(_04398_));
 sky130_fd_sc_hd__a2111oi_2 _09692_ (.A1(_04393_),
    .A2(_04394_),
    .B1(_03825_),
    .C1(_04396_),
    .D1(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__clkinv_1 _09699_ (.A(net595),
    .Y(_04406_));
 sky130_fd_sc_hd__mux2i_1 _09702_ (.A0(\core.CPU_Xreg_value_a4[11][0] ),
    .A1(\core.CPU_Xreg_value_a4[27][0] ),
    .S(\core.CPU_rf_rd_index1_a2[4] ),
    .Y(_04409_));
 sky130_fd_sc_hd__inv_1 _09703_ (.A(\core.CPU_rf_rd_index1_a2[4] ),
    .Y(_04410_));
 sky130_fd_sc_hd__nor2_1 _09704_ (.A(net596),
    .B(net543),
    .Y(_04411_));
 sky130_fd_sc_hd__nand2_1 _09705_ (.A(net620),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__o21ai_0 _09706_ (.A1(net544),
    .A2(_04409_),
    .B1(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__mux2_2 _09708_ (.A0(\core.CPU_Xreg_value_a4[10][0] ),
    .A1(\core.CPU_Xreg_value_a4[26][0] ),
    .S(net593),
    .X(_04415_));
 sky130_fd_sc_hd__nor2_1 _09709_ (.A(net545),
    .B(\core.CPU_rf_rd_index1_a2[0] ),
    .Y(_04416_));
 sky130_fd_sc_hd__clkinv_1 _09712_ (.A(\core.CPU_rf_rd_index1_a2[0] ),
    .Y(_04419_));
 sky130_fd_sc_hd__inv_1 _09715_ (.A(\core.CPU_Xreg_value_a4[1][0] ),
    .Y(_04422_));
 sky130_fd_sc_hd__a21oi_1 _09717_ (.A1(net598),
    .A2(_04422_),
    .B1(net593),
    .Y(_04424_));
 sky130_fd_sc_hd__a21oi_1 _09718_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[16][0] ),
    .B1(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__nor2_1 _09719_ (.A(net596),
    .B(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__a221oi_1 _09720_ (.A1(net598),
    .A2(_04413_),
    .B1(_04415_),
    .B2(net471),
    .C1(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__nor2_1 _09721_ (.A(net596),
    .B(net593),
    .Y(_04428_));
 sky130_fd_sc_hd__nand2_1 _09722_ (.A(net542),
    .B(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__nor2_1 _09724_ (.A(\core.CPU_Xreg_value_a4[0][0] ),
    .B(net469),
    .Y(_04431_));
 sky130_fd_sc_hd__nor2_1 _09725_ (.A(_04427_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__nor2_1 _09726_ (.A(net434),
    .B(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__a21oi_1 _09727_ (.A1(net394),
    .A2(net434),
    .B1(_04433_),
    .Y(\core.CPU_src1_value_a2[0] ));
 sky130_fd_sc_hd__mux2_2 _09729_ (.A0(\core.CPU_Xreg_value_a4[16][10] ),
    .A1(\core.CPU_Xreg_value_a4[17][10] ),
    .S(net598),
    .X(_04435_));
 sky130_fd_sc_hd__nor2_1 _09730_ (.A(\core.CPU_rf_rd_index1_a2[4] ),
    .B(net598),
    .Y(_04436_));
 sky130_fd_sc_hd__a221oi_1 _09731_ (.A1(\core.CPU_rf_rd_index1_a2[4] ),
    .A2(_04435_),
    .B1(_04436_),
    .B2(\core.CPU_Xreg_value_a4[0][10] ),
    .C1(net596),
    .Y(_04437_));
 sky130_fd_sc_hd__mux2_2 _09732_ (.A0(\core.CPU_Xreg_value_a4[26][10] ),
    .A1(\core.CPU_Xreg_value_a4[27][10] ),
    .S(net598),
    .X(_04438_));
 sky130_fd_sc_hd__nor2_2 _09733_ (.A(\core.CPU_rf_rd_index1_a2[4] ),
    .B(net542),
    .Y(_04439_));
 sky130_fd_sc_hd__a221oi_1 _09735_ (.A1(\core.CPU_rf_rd_index1_a2[4] ),
    .A2(_04438_),
    .B1(net468),
    .B2(\core.CPU_Xreg_value_a4[11][10] ),
    .C1(net544),
    .Y(_04441_));
 sky130_fd_sc_hd__nor2_2 _09736_ (.A(net596),
    .B(net542),
    .Y(_04442_));
 sky130_fd_sc_hd__a22oi_1 _09737_ (.A1(\core.CPU_Xreg_value_a4[10][10] ),
    .A2(net471),
    .B1(_04442_),
    .B2(\core.CPU_Xreg_value_a4[1][10] ),
    .Y(_04443_));
 sky130_fd_sc_hd__o22ai_1 _09739_ (.A1(_04437_),
    .A2(_04441_),
    .B1(_04443_),
    .B2(\core.CPU_rf_rd_index1_a2[4] ),
    .Y(_04445_));
 sky130_fd_sc_hd__nor2_1 _09740_ (.A(net432),
    .B(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__a21oi_1 _09741_ (.A1(_02640_),
    .A2(net432),
    .B1(_04446_),
    .Y(\core.CPU_src1_value_a2[10] ));
 sky130_fd_sc_hd__nand2_1 _09746_ (.A(net543),
    .B(net598),
    .Y(_04451_));
 sky130_fd_sc_hd__mux2_2 _09747_ (.A0(\core.CPU_Xreg_value_a4[16][11] ),
    .A1(\core.CPU_Xreg_value_a4[17][11] ),
    .S(net598),
    .X(_04452_));
 sky130_fd_sc_hd__o22ai_1 _09750_ (.A1(\core.CPU_Xreg_value_a4[1][11] ),
    .A2(_04451_),
    .B1(_04452_),
    .B2(net543),
    .Y(_04455_));
 sky130_fd_sc_hd__mux4_2 _09752_ (.A0(\core.CPU_Xreg_value_a4[10][11] ),
    .A1(\core.CPU_Xreg_value_a4[11][11] ),
    .A2(\core.CPU_Xreg_value_a4[26][11] ),
    .A3(\core.CPU_Xreg_value_a4[27][11] ),
    .S0(net598),
    .S1(\core.CPU_rf_rd_index1_a2[4] ),
    .X(_04457_));
 sky130_fd_sc_hd__nor2_1 _09753_ (.A(net544),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__a21oi_1 _09754_ (.A1(net544),
    .A2(_04455_),
    .B1(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__o21ai_1 _09755_ (.A1(\core.CPU_Xreg_value_a4[0][11] ),
    .A2(net469),
    .B1(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__nand2_1 _09757_ (.A(_02717_),
    .B(net432),
    .Y(_04462_));
 sky130_fd_sc_hd__o21ai_0 _09758_ (.A1(net432),
    .A2(net408),
    .B1(_04462_),
    .Y(\core.CPU_src1_value_a2[11] ));
 sky130_fd_sc_hd__o21ai_0 _09760_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[1][12] ),
    .B1(net543),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2_1 _09762_ (.A(net542),
    .B(\core.CPU_Xreg_value_a4[16][12] ),
    .Y(_04466_));
 sky130_fd_sc_hd__a21oi_1 _09763_ (.A1(_04464_),
    .A2(_04466_),
    .B1(net595),
    .Y(_04467_));
 sky130_fd_sc_hd__mux2_2 _09765_ (.A0(\core.CPU_Xreg_value_a4[11][12] ),
    .A1(\core.CPU_Xreg_value_a4[27][12] ),
    .S(net593),
    .X(_04469_));
 sky130_fd_sc_hd__a221oi_1 _09767_ (.A1(\core.CPU_Xreg_value_a4[17][12] ),
    .A2(net472),
    .B1(_04469_),
    .B2(net595),
    .C1(net542),
    .Y(_04471_));
 sky130_fd_sc_hd__nor2_1 _09768_ (.A(net545),
    .B(net543),
    .Y(_04472_));
 sky130_fd_sc_hd__a221oi_1 _09769_ (.A1(net543),
    .A2(\core.CPU_Xreg_value_a4[10][12] ),
    .B1(net466),
    .B2(\core.CPU_Xreg_value_a4[26][12] ),
    .C1(net597),
    .Y(_04473_));
 sky130_fd_sc_hd__nor2_1 _09770_ (.A(_04471_),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__o22ai_1 _09771_ (.A1(\core.CPU_Xreg_value_a4[0][12] ),
    .A2(net470),
    .B1(_04467_),
    .B2(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__a21boi_0 _09772_ (.A1(net611),
    .A2(_02763_),
    .B1_N(net370),
    .Y(_04476_));
 sky130_fd_sc_hd__mux2i_1 _09774_ (.A0(_04475_),
    .A1(_04476_),
    .S(net432),
    .Y(\core.CPU_src1_value_a2[12] ));
 sky130_fd_sc_hd__mux2_2 _09775_ (.A0(\core.CPU_Xreg_value_a4[0][13] ),
    .A1(\core.CPU_Xreg_value_a4[16][13] ),
    .S(net594),
    .X(_04478_));
 sky130_fd_sc_hd__nor2_1 _09776_ (.A(net595),
    .B(\core.CPU_rf_rd_index1_a2[0] ),
    .Y(_04479_));
 sky130_fd_sc_hd__mux2_2 _09777_ (.A0(\core.CPU_Xreg_value_a4[26][13] ),
    .A1(\core.CPU_Xreg_value_a4[27][13] ),
    .S(net597),
    .X(_04480_));
 sky130_fd_sc_hd__a22oi_1 _09779_ (.A1(\core.CPU_Xreg_value_a4[10][13] ),
    .A2(net541),
    .B1(_04480_),
    .B2(net594),
    .Y(_04482_));
 sky130_fd_sc_hd__nor2_1 _09780_ (.A(net545),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__nor2_1 _09781_ (.A(net545),
    .B(net593),
    .Y(_04484_));
 sky130_fd_sc_hd__mux2i_1 _09783_ (.A0(\core.CPU_Xreg_value_a4[1][13] ),
    .A1(\core.CPU_Xreg_value_a4[17][13] ),
    .S(net594),
    .Y(_04486_));
 sky130_fd_sc_hd__nor2_1 _09784_ (.A(net595),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__a21oi_1 _09785_ (.A1(\core.CPU_Xreg_value_a4[11][13] ),
    .A2(_04484_),
    .B1(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__nor2_1 _09786_ (.A(_04419_),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__a2111oi_0 _09787_ (.A1(_04478_),
    .A2(_04479_),
    .B1(_04483_),
    .C1(_04489_),
    .D1(net432),
    .Y(_04490_));
 sky130_fd_sc_hd__a21oi_1 _09788_ (.A1(_02810_),
    .A2(net433),
    .B1(net407),
    .Y(\core.CPU_src1_value_a2[13] ));
 sky130_fd_sc_hd__nand2_1 _09790_ (.A(net544),
    .B(net598),
    .Y(_04492_));
 sky130_fd_sc_hd__mux2_2 _09791_ (.A0(\core.CPU_Xreg_value_a4[10][14] ),
    .A1(\core.CPU_Xreg_value_a4[11][14] ),
    .S(net598),
    .X(_04493_));
 sky130_fd_sc_hd__o22ai_1 _09792_ (.A1(\core.CPU_Xreg_value_a4[1][14] ),
    .A2(net465),
    .B1(_04493_),
    .B2(net544),
    .Y(_04494_));
 sky130_fd_sc_hd__mux4_2 _09793_ (.A0(\core.CPU_Xreg_value_a4[16][14] ),
    .A1(\core.CPU_Xreg_value_a4[17][14] ),
    .A2(\core.CPU_Xreg_value_a4[26][14] ),
    .A3(\core.CPU_Xreg_value_a4[27][14] ),
    .S0(net598),
    .S1(net596),
    .X(_04495_));
 sky130_fd_sc_hd__nor2_1 _09794_ (.A(net543),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__a21oi_1 _09795_ (.A1(net543),
    .A2(_04494_),
    .B1(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__o21ai_2 _09796_ (.A1(\core.CPU_Xreg_value_a4[0][14] ),
    .A2(net469),
    .B1(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__mux2i_1 _09797_ (.A0(net406),
    .A1(_02866_),
    .S(net432),
    .Y(\core.CPU_src1_value_a2[14] ));
 sky130_fd_sc_hd__o21ai_0 _09798_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[1][15] ),
    .B1(net543),
    .Y(_04499_));
 sky130_fd_sc_hd__nand2_1 _09799_ (.A(net542),
    .B(\core.CPU_Xreg_value_a4[16][15] ),
    .Y(_04500_));
 sky130_fd_sc_hd__a21oi_1 _09800_ (.A1(_04499_),
    .A2(_04500_),
    .B1(net595),
    .Y(_04501_));
 sky130_fd_sc_hd__mux2_2 _09801_ (.A0(\core.CPU_Xreg_value_a4[11][15] ),
    .A1(\core.CPU_Xreg_value_a4[27][15] ),
    .S(net593),
    .X(_04502_));
 sky130_fd_sc_hd__a221oi_1 _09802_ (.A1(\core.CPU_Xreg_value_a4[17][15] ),
    .A2(net472),
    .B1(_04502_),
    .B2(net595),
    .C1(net542),
    .Y(_04503_));
 sky130_fd_sc_hd__a221oi_1 _09803_ (.A1(net543),
    .A2(\core.CPU_Xreg_value_a4[10][15] ),
    .B1(net466),
    .B2(\core.CPU_Xreg_value_a4[26][15] ),
    .C1(\core.CPU_rf_rd_index1_a2[0] ),
    .Y(_04504_));
 sky130_fd_sc_hd__nor2_1 _09804_ (.A(_04503_),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__o22ai_1 _09805_ (.A1(\core.CPU_Xreg_value_a4[0][15] ),
    .A2(net470),
    .B1(_04501_),
    .B2(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__mux2i_1 _09806_ (.A0(_04506_),
    .A1(_02909_),
    .S(net433),
    .Y(\core.CPU_src1_value_a2[15] ));
 sky130_fd_sc_hd__a22oi_1 _09807_ (.A1(\core.CPU_Xreg_value_a4[0][16] ),
    .A2(_04428_),
    .B1(net466),
    .B2(\core.CPU_Xreg_value_a4[26][16] ),
    .Y(_04507_));
 sky130_fd_sc_hd__mux2_2 _09808_ (.A0(\core.CPU_Xreg_value_a4[16][16] ),
    .A1(\core.CPU_Xreg_value_a4[17][16] ),
    .S(net597),
    .X(_04508_));
 sky130_fd_sc_hd__mux2i_1 _09809_ (.A0(\core.CPU_Xreg_value_a4[11][16] ),
    .A1(\core.CPU_Xreg_value_a4[27][16] ),
    .S(net593),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_1 _09810_ (.A(net595),
    .B(net597),
    .Y(_04510_));
 sky130_fd_sc_hd__a22oi_1 _09811_ (.A1(\core.CPU_Xreg_value_a4[10][16] ),
    .A2(net471),
    .B1(net467),
    .B2(\core.CPU_Xreg_value_a4[1][16] ),
    .Y(_04511_));
 sky130_fd_sc_hd__o22ai_1 _09812_ (.A1(_04509_),
    .A2(_04510_),
    .B1(_04511_),
    .B2(net593),
    .Y(_04512_));
 sky130_fd_sc_hd__a21oi_1 _09813_ (.A1(net472),
    .A2(_04508_),
    .B1(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__o21ai_0 _09814_ (.A1(net597),
    .A2(_04507_),
    .B1(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__mux2_2 _09815_ (.A0(net388),
    .A1(_02956_),
    .S(net433),
    .X(\core.CPU_src1_value_a2[16] ));
 sky130_fd_sc_hd__mux2i_1 _09816_ (.A0(\core.CPU_Xreg_value_a4[11][17] ),
    .A1(\core.CPU_Xreg_value_a4[27][17] ),
    .S(net594),
    .Y(_04515_));
 sky130_fd_sc_hd__nand2_1 _09817_ (.A(\core.CPU_Xreg_value_a4[17][17] ),
    .B(net472),
    .Y(_04516_));
 sky130_fd_sc_hd__o21ai_0 _09818_ (.A1(net545),
    .A2(_04515_),
    .B1(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__o21ai_0 _09819_ (.A1(_04419_),
    .A2(\core.CPU_Xreg_value_a4[1][17] ),
    .B1(net545),
    .Y(_04518_));
 sky130_fd_sc_hd__a21boi_0 _09820_ (.A1(_04419_),
    .A2(\core.CPU_Xreg_value_a4[10][17] ),
    .B1_N(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__mux2i_1 _09821_ (.A0(\core.CPU_Xreg_value_a4[16][17] ),
    .A1(\core.CPU_Xreg_value_a4[26][17] ),
    .S(net595),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _09822_ (.A(\core.CPU_rf_rd_index1_a2[4] ),
    .B(net542),
    .Y(_04521_));
 sky130_fd_sc_hd__o22ai_1 _09823_ (.A1(net594),
    .A2(_04519_),
    .B1(_04520_),
    .B2(net464),
    .Y(_04522_));
 sky130_fd_sc_hd__a21oi_1 _09824_ (.A1(net597),
    .A2(_04517_),
    .B1(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__nor2_1 _09825_ (.A(\core.CPU_Xreg_value_a4[0][17] ),
    .B(net470),
    .Y(_04524_));
 sky130_fd_sc_hd__nor2_1 _09826_ (.A(_04523_),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__nor2_1 _09827_ (.A(net433),
    .B(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__a21oi_1 _09828_ (.A1(_03003_),
    .A2(net433),
    .B1(_04526_),
    .Y(\core.CPU_src1_value_a2[17] ));
 sky130_fd_sc_hd__mux2_2 _09829_ (.A0(\core.CPU_Xreg_value_a4[0][18] ),
    .A1(\core.CPU_Xreg_value_a4[16][18] ),
    .S(net594),
    .X(_04527_));
 sky130_fd_sc_hd__a221oi_1 _09830_ (.A1(\core.CPU_Xreg_value_a4[10][18] ),
    .A2(net471),
    .B1(net467),
    .B2(\core.CPU_Xreg_value_a4[1][18] ),
    .C1(net594),
    .Y(_04528_));
 sky130_fd_sc_hd__a221oi_1 _09831_ (.A1(\core.CPU_Xreg_value_a4[26][18] ),
    .A2(net471),
    .B1(net467),
    .B2(\core.CPU_Xreg_value_a4[17][18] ),
    .C1(net543),
    .Y(_04529_));
 sky130_fd_sc_hd__nor2_1 _09832_ (.A(_04528_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__mux2i_1 _09833_ (.A0(\core.CPU_Xreg_value_a4[11][18] ),
    .A1(\core.CPU_Xreg_value_a4[27][18] ),
    .S(net594),
    .Y(_04531_));
 sky130_fd_sc_hd__nor2_1 _09834_ (.A(_04510_),
    .B(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__a2111oi_0 _09835_ (.A1(_04479_),
    .A2(_04527_),
    .B1(_04530_),
    .C1(net432),
    .D1(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__a21oi_1 _09836_ (.A1(net359),
    .A2(net433),
    .B1(net405),
    .Y(\core.CPU_src1_value_a2[18] ));
 sky130_fd_sc_hd__a21o_1 _09837_ (.A1(net476),
    .A2(_03055_),
    .B1(_03089_),
    .X(_04534_));
 sky130_fd_sc_hd__mux2i_1 _09838_ (.A0(\core.CPU_Xreg_value_a4[11][19] ),
    .A1(\core.CPU_Xreg_value_a4[27][19] ),
    .S(net594),
    .Y(_04535_));
 sky130_fd_sc_hd__nand2_1 _09839_ (.A(\core.CPU_Xreg_value_a4[17][19] ),
    .B(net472),
    .Y(_04536_));
 sky130_fd_sc_hd__o21ai_0 _09840_ (.A1(net545),
    .A2(_04535_),
    .B1(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__o21ai_0 _09841_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[1][19] ),
    .B1(net545),
    .Y(_04538_));
 sky130_fd_sc_hd__a21boi_0 _09842_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[10][19] ),
    .B1_N(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__mux2i_1 _09843_ (.A0(\core.CPU_Xreg_value_a4[16][19] ),
    .A1(\core.CPU_Xreg_value_a4[26][19] ),
    .S(net595),
    .Y(_04540_));
 sky130_fd_sc_hd__o22ai_1 _09844_ (.A1(net593),
    .A2(_04539_),
    .B1(_04540_),
    .B2(net464),
    .Y(_04541_));
 sky130_fd_sc_hd__a21oi_1 _09845_ (.A1(\core.CPU_rf_rd_index1_a2[0] ),
    .A2(_04537_),
    .B1(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__nor2_1 _09846_ (.A(\core.CPU_Xreg_value_a4[0][19] ),
    .B(net470),
    .Y(_04543_));
 sky130_fd_sc_hd__nor2_1 _09847_ (.A(_04542_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__nor2_1 _09848_ (.A(net432),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__a21oi_1 _09849_ (.A1(net432),
    .A2(_04534_),
    .B1(_04545_),
    .Y(\core.CPU_src1_value_a2[19] ));
 sky130_fd_sc_hd__o21ai_0 _09850_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[1][1] ),
    .B1(net543),
    .Y(_04546_));
 sky130_fd_sc_hd__nand2_1 _09851_ (.A(net542),
    .B(\core.CPU_Xreg_value_a4[16][1] ),
    .Y(_04547_));
 sky130_fd_sc_hd__a21oi_1 _09852_ (.A1(_04546_),
    .A2(_04547_),
    .B1(net596),
    .Y(_04548_));
 sky130_fd_sc_hd__mux2_2 _09853_ (.A0(\core.CPU_Xreg_value_a4[11][1] ),
    .A1(\core.CPU_Xreg_value_a4[27][1] ),
    .S(net593),
    .X(_04549_));
 sky130_fd_sc_hd__a221oi_1 _09854_ (.A1(\core.CPU_Xreg_value_a4[17][1] ),
    .A2(net472),
    .B1(_04549_),
    .B2(net596),
    .C1(net542),
    .Y(_04550_));
 sky130_fd_sc_hd__a221oi_1 _09855_ (.A1(net543),
    .A2(\core.CPU_Xreg_value_a4[10][1] ),
    .B1(_04472_),
    .B2(\core.CPU_Xreg_value_a4[26][1] ),
    .C1(\core.CPU_rf_rd_index1_a2[0] ),
    .Y(_04551_));
 sky130_fd_sc_hd__nor2_1 _09856_ (.A(_04550_),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__o22ai_1 _09857_ (.A1(\core.CPU_Xreg_value_a4[0][1] ),
    .A2(net469),
    .B1(_04548_),
    .B2(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__nand2_1 _09858_ (.A(_03099_),
    .B(net432),
    .Y(_04554_));
 sky130_fd_sc_hd__o21ai_0 _09859_ (.A1(net432),
    .A2(net404),
    .B1(_04554_),
    .Y(\core.CPU_src1_value_a2[1] ));
 sky130_fd_sc_hd__mux2_2 _09860_ (.A0(\core.CPU_Xreg_value_a4[10][20] ),
    .A1(\core.CPU_Xreg_value_a4[11][20] ),
    .S(net598),
    .X(_04555_));
 sky130_fd_sc_hd__o22ai_1 _09861_ (.A1(\core.CPU_Xreg_value_a4[1][20] ),
    .A2(net465),
    .B1(_04555_),
    .B2(net544),
    .Y(_04556_));
 sky130_fd_sc_hd__mux4_2 _09862_ (.A0(\core.CPU_Xreg_value_a4[16][20] ),
    .A1(\core.CPU_Xreg_value_a4[17][20] ),
    .A2(\core.CPU_Xreg_value_a4[26][20] ),
    .A3(\core.CPU_Xreg_value_a4[27][20] ),
    .S0(net598),
    .S1(net596),
    .X(_04557_));
 sky130_fd_sc_hd__nor2_1 _09863_ (.A(net543),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__a21oi_1 _09864_ (.A1(net543),
    .A2(_04556_),
    .B1(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__o21ai_1 _09865_ (.A1(\core.CPU_Xreg_value_a4[0][20] ),
    .A2(net469),
    .B1(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__nand2_1 _09866_ (.A(_03141_),
    .B(net432),
    .Y(_04561_));
 sky130_fd_sc_hd__o21ai_0 _09867_ (.A1(net432),
    .A2(net403),
    .B1(_04561_),
    .Y(\core.CPU_src1_value_a2[20] ));
 sky130_fd_sc_hd__o21ai_0 _09868_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[1][21] ),
    .B1(net544),
    .Y(_04562_));
 sky130_fd_sc_hd__a21boi_0 _09869_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[10][21] ),
    .B1_N(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__mux2i_1 _09870_ (.A0(\core.CPU_Xreg_value_a4[16][21] ),
    .A1(\core.CPU_Xreg_value_a4[26][21] ),
    .S(net596),
    .Y(_04564_));
 sky130_fd_sc_hd__mux2i_1 _09871_ (.A0(\core.CPU_Xreg_value_a4[11][21] ),
    .A1(\core.CPU_Xreg_value_a4[27][21] ),
    .S(\core.CPU_rf_rd_index1_a2[4] ),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _09872_ (.A(\core.CPU_Xreg_value_a4[17][21] ),
    .B(_04411_),
    .Y(_04566_));
 sky130_fd_sc_hd__o21ai_0 _09873_ (.A1(net544),
    .A2(_04565_),
    .B1(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__nand2_1 _09874_ (.A(net598),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__o221ai_1 _09875_ (.A1(\core.CPU_rf_rd_index1_a2[4] ),
    .A2(_04563_),
    .B1(_04564_),
    .B2(_04521_),
    .C1(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__o21ai_1 _09876_ (.A1(\core.CPU_Xreg_value_a4[0][21] ),
    .A2(net469),
    .B1(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__nand2_1 _09877_ (.A(_03188_),
    .B(net432),
    .Y(_04571_));
 sky130_fd_sc_hd__o21ai_0 _09878_ (.A1(net432),
    .A2(net381),
    .B1(_04571_),
    .Y(\core.CPU_src1_value_a2[21] ));
 sky130_fd_sc_hd__mux2_2 _09879_ (.A0(\core.CPU_Xreg_value_a4[16][22] ),
    .A1(\core.CPU_Xreg_value_a4[17][22] ),
    .S(\core.CPU_rf_rd_index1_a2[0] ),
    .X(_04572_));
 sky130_fd_sc_hd__o22ai_1 _09880_ (.A1(\core.CPU_Xreg_value_a4[1][22] ),
    .A2(_04451_),
    .B1(_04572_),
    .B2(net543),
    .Y(_04573_));
 sky130_fd_sc_hd__mux4_2 _09881_ (.A0(\core.CPU_Xreg_value_a4[10][22] ),
    .A1(\core.CPU_Xreg_value_a4[11][22] ),
    .A2(\core.CPU_Xreg_value_a4[26][22] ),
    .A3(\core.CPU_Xreg_value_a4[27][22] ),
    .S0(\core.CPU_rf_rd_index1_a2[0] ),
    .S1(net593),
    .X(_04574_));
 sky130_fd_sc_hd__nor2_1 _09882_ (.A(net545),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21oi_1 _09883_ (.A1(net545),
    .A2(_04573_),
    .B1(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__o21ai_0 _09884_ (.A1(\core.CPU_Xreg_value_a4[0][22] ),
    .A2(net470),
    .B1(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__and2_1 _09885_ (.A(_03211_),
    .B(net369),
    .X(_04578_));
 sky130_fd_sc_hd__mux2i_1 _09886_ (.A0(_04577_),
    .A1(_04578_),
    .S(net433),
    .Y(\core.CPU_src1_value_a2[22] ));
 sky130_fd_sc_hd__and2_1 _09887_ (.A(_03241_),
    .B(_03274_),
    .X(_04579_));
 sky130_fd_sc_hd__mux2_2 _09888_ (.A0(\core.CPU_Xreg_value_a4[0][23] ),
    .A1(\core.CPU_Xreg_value_a4[16][23] ),
    .S(net594),
    .X(_04580_));
 sky130_fd_sc_hd__mux2_2 _09889_ (.A0(\core.CPU_Xreg_value_a4[26][23] ),
    .A1(\core.CPU_Xreg_value_a4[27][23] ),
    .S(net597),
    .X(_04581_));
 sky130_fd_sc_hd__a22oi_1 _09890_ (.A1(\core.CPU_Xreg_value_a4[10][23] ),
    .A2(net541),
    .B1(_04581_),
    .B2(net594),
    .Y(_04582_));
 sky130_fd_sc_hd__nor2_1 _09891_ (.A(net545),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__mux2i_1 _09892_ (.A0(\core.CPU_Xreg_value_a4[1][23] ),
    .A1(\core.CPU_Xreg_value_a4[17][23] ),
    .S(net594),
    .Y(_04584_));
 sky130_fd_sc_hd__nor2_1 _09893_ (.A(net595),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__a21oi_1 _09894_ (.A1(\core.CPU_Xreg_value_a4[11][23] ),
    .A2(_04484_),
    .B1(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__nor2_1 _09895_ (.A(_04419_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__a2111oi_0 _09896_ (.A1(_04479_),
    .A2(_04580_),
    .B1(_04583_),
    .C1(_04587_),
    .D1(net432),
    .Y(_04588_));
 sky130_fd_sc_hd__a21oi_1 _09897_ (.A1(_04579_),
    .A2(net433),
    .B1(net402),
    .Y(\core.CPU_src1_value_a2[23] ));
 sky130_fd_sc_hd__a21boi_0 _09898_ (.A1(net476),
    .A2(_03307_),
    .B1_N(_03301_),
    .Y(_04589_));
 sky130_fd_sc_hd__mux2i_1 _09899_ (.A0(\core.CPU_Xreg_value_a4[11][24] ),
    .A1(\core.CPU_Xreg_value_a4[27][24] ),
    .S(net594),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_1 _09900_ (.A(\core.CPU_Xreg_value_a4[17][24] ),
    .B(net472),
    .Y(_04591_));
 sky130_fd_sc_hd__o21ai_0 _09901_ (.A1(net545),
    .A2(_04590_),
    .B1(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__o21ai_0 _09902_ (.A1(_04419_),
    .A2(\core.CPU_Xreg_value_a4[1][24] ),
    .B1(net545),
    .Y(_04593_));
 sky130_fd_sc_hd__a21boi_0 _09903_ (.A1(_04419_),
    .A2(\core.CPU_Xreg_value_a4[10][24] ),
    .B1_N(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__mux2i_1 _09904_ (.A0(\core.CPU_Xreg_value_a4[16][24] ),
    .A1(\core.CPU_Xreg_value_a4[26][24] ),
    .S(net595),
    .Y(_04595_));
 sky130_fd_sc_hd__o22ai_1 _09905_ (.A1(net594),
    .A2(_04594_),
    .B1(_04595_),
    .B2(net464),
    .Y(_04596_));
 sky130_fd_sc_hd__a21oi_1 _09906_ (.A1(net597),
    .A2(_04592_),
    .B1(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__nor2_1 _09907_ (.A(\core.CPU_Xreg_value_a4[0][24] ),
    .B(net470),
    .Y(_04598_));
 sky130_fd_sc_hd__nor3_1 _09908_ (.A(net432),
    .B(_04597_),
    .C(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__a21o_1 _09909_ (.A1(_04589_),
    .A2(net433),
    .B1(_04599_),
    .X(\core.CPU_src1_value_a2[24] ));
 sky130_fd_sc_hd__o21ai_0 _09910_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[1][25] ),
    .B1(net543),
    .Y(_04600_));
 sky130_fd_sc_hd__nand2_1 _09911_ (.A(net542),
    .B(\core.CPU_Xreg_value_a4[16][25] ),
    .Y(_04601_));
 sky130_fd_sc_hd__a21oi_1 _09912_ (.A1(_04600_),
    .A2(_04601_),
    .B1(net595),
    .Y(_04602_));
 sky130_fd_sc_hd__mux2_2 _09913_ (.A0(\core.CPU_Xreg_value_a4[11][25] ),
    .A1(\core.CPU_Xreg_value_a4[27][25] ),
    .S(net593),
    .X(_04603_));
 sky130_fd_sc_hd__a221oi_1 _09914_ (.A1(\core.CPU_Xreg_value_a4[17][25] ),
    .A2(net472),
    .B1(_04603_),
    .B2(net595),
    .C1(net542),
    .Y(_04604_));
 sky130_fd_sc_hd__a221oi_1 _09915_ (.A1(net543),
    .A2(\core.CPU_Xreg_value_a4[10][25] ),
    .B1(net466),
    .B2(\core.CPU_Xreg_value_a4[26][25] ),
    .C1(\core.CPU_rf_rd_index1_a2[0] ),
    .Y(_04605_));
 sky130_fd_sc_hd__nor2_1 _09916_ (.A(_04604_),
    .B(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__o22ai_1 _09917_ (.A1(\core.CPU_Xreg_value_a4[0][25] ),
    .A2(net469),
    .B1(_04602_),
    .B2(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__nand2_1 _09918_ (.A(_03352_),
    .B(net433),
    .Y(_04608_));
 sky130_fd_sc_hd__o21ai_0 _09919_ (.A1(net433),
    .A2(_04607_),
    .B1(_04608_),
    .Y(\core.CPU_src1_value_a2[25] ));
 sky130_fd_sc_hd__mux4_2 _09920_ (.A0(\core.CPU_Xreg_value_a4[16][26] ),
    .A1(\core.CPU_Xreg_value_a4[17][26] ),
    .A2(\core.CPU_Xreg_value_a4[26][26] ),
    .A3(\core.CPU_Xreg_value_a4[27][26] ),
    .S0(net597),
    .S1(net595),
    .X(_04609_));
 sky130_fd_sc_hd__inv_1 _09921_ (.A(\core.CPU_Xreg_value_a4[1][26] ),
    .Y(_04610_));
 sky130_fd_sc_hd__mux2i_1 _09922_ (.A0(\core.CPU_Xreg_value_a4[10][26] ),
    .A1(\core.CPU_Xreg_value_a4[11][26] ),
    .S(net597),
    .Y(_04611_));
 sky130_fd_sc_hd__a221oi_1 _09923_ (.A1(_04610_),
    .A2(net467),
    .B1(_04611_),
    .B2(net595),
    .C1(net594),
    .Y(_04612_));
 sky130_fd_sc_hd__a21oi_1 _09924_ (.A1(net594),
    .A2(_04609_),
    .B1(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__nor2_1 _09925_ (.A(\core.CPU_Xreg_value_a4[0][26] ),
    .B(net470),
    .Y(_04614_));
 sky130_fd_sc_hd__nor2_1 _09926_ (.A(_04613_),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__nor2_1 _09927_ (.A(net433),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__a21oi_1 _09928_ (.A1(_03387_),
    .A2(net433),
    .B1(_04616_),
    .Y(\core.CPU_src1_value_a2[26] ));
 sky130_fd_sc_hd__mux4_2 _09929_ (.A0(\core.CPU_Xreg_value_a4[16][27] ),
    .A1(\core.CPU_Xreg_value_a4[17][27] ),
    .A2(\core.CPU_Xreg_value_a4[26][27] ),
    .A3(\core.CPU_Xreg_value_a4[27][27] ),
    .S0(net597),
    .S1(net595),
    .X(_04617_));
 sky130_fd_sc_hd__nand2_1 _09930_ (.A(net594),
    .B(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__mux2_2 _09931_ (.A0(\core.CPU_Xreg_value_a4[10][27] ),
    .A1(\core.CPU_Xreg_value_a4[11][27] ),
    .S(net597),
    .X(_04619_));
 sky130_fd_sc_hd__o221ai_1 _09932_ (.A1(\core.CPU_Xreg_value_a4[1][27] ),
    .A2(net465),
    .B1(_04619_),
    .B2(net545),
    .C1(net543),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _09933_ (.A(\core.CPU_Xreg_value_a4[0][27] ),
    .B(net470),
    .Y(_04621_));
 sky130_fd_sc_hd__a21oi_1 _09934_ (.A1(_04618_),
    .A2(_04620_),
    .B1(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__nor2_1 _09935_ (.A(net433),
    .B(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__a31oi_1 _09936_ (.A1(net353),
    .A2(_03431_),
    .A3(net433),
    .B1(_04623_),
    .Y(\core.CPU_src1_value_a2[27] ));
 sky130_fd_sc_hd__nand2_1 _09937_ (.A(_02794_),
    .B(_03462_),
    .Y(_04624_));
 sky130_fd_sc_hd__a21oi_1 _09938_ (.A1(net557),
    .A2(_03457_),
    .B1(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__o21ai_0 _09939_ (.A1(_03457_),
    .A2(net391),
    .B1(net433),
    .Y(_04626_));
 sky130_fd_sc_hd__inv_1 _09940_ (.A(\core.CPU_Xreg_value_a4[26][28] ),
    .Y(_04627_));
 sky130_fd_sc_hd__nand2_1 _09941_ (.A(\core.CPU_Xreg_value_a4[11][28] ),
    .B(net468),
    .Y(_04628_));
 sky130_fd_sc_hd__o21ai_0 _09942_ (.A1(_04627_),
    .A2(net464),
    .B1(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__nand2_1 _09943_ (.A(net595),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__inv_1 _09944_ (.A(\core.CPU_Xreg_value_a4[10][28] ),
    .Y(_04631_));
 sky130_fd_sc_hd__o21ai_0 _09945_ (.A1(_04419_),
    .A2(\core.CPU_Xreg_value_a4[1][28] ),
    .B1(net545),
    .Y(_04632_));
 sky130_fd_sc_hd__o21ai_0 _09946_ (.A1(net597),
    .A2(_04631_),
    .B1(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__mux2i_1 _09947_ (.A0(\core.CPU_Xreg_value_a4[16][28] ),
    .A1(\core.CPU_Xreg_value_a4[17][28] ),
    .S(net597),
    .Y(_04634_));
 sky130_fd_sc_hd__nand3_1 _09948_ (.A(net595),
    .B(net597),
    .C(\core.CPU_Xreg_value_a4[27][28] ),
    .Y(_04635_));
 sky130_fd_sc_hd__o211ai_1 _09949_ (.A1(net595),
    .A2(_04634_),
    .B1(_04635_),
    .C1(net594),
    .Y(_04636_));
 sky130_fd_sc_hd__o21ai_0 _09950_ (.A1(net594),
    .A2(_04633_),
    .B1(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__nor2_1 _09951_ (.A(\core.CPU_Xreg_value_a4[0][28] ),
    .B(net470),
    .Y(_04638_));
 sky130_fd_sc_hd__a21oi_1 _09952_ (.A1(_04630_),
    .A2(_04637_),
    .B1(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__o22a_1 _09953_ (.A1(_04625_),
    .A2(_04626_),
    .B1(_04639_),
    .B2(net433),
    .X(\core.CPU_src1_value_a2[28] ));
 sky130_fd_sc_hd__mux2_2 _09954_ (.A0(\core.CPU_Xreg_value_a4[10][29] ),
    .A1(\core.CPU_Xreg_value_a4[11][29] ),
    .S(net598),
    .X(_04640_));
 sky130_fd_sc_hd__o22ai_1 _09955_ (.A1(\core.CPU_Xreg_value_a4[1][29] ),
    .A2(net465),
    .B1(_04640_),
    .B2(net544),
    .Y(_04641_));
 sky130_fd_sc_hd__mux4_2 _09956_ (.A0(\core.CPU_Xreg_value_a4[16][29] ),
    .A1(\core.CPU_Xreg_value_a4[17][29] ),
    .A2(\core.CPU_Xreg_value_a4[26][29] ),
    .A3(\core.CPU_Xreg_value_a4[27][29] ),
    .S0(net598),
    .S1(net596),
    .X(_04642_));
 sky130_fd_sc_hd__nor2_1 _09957_ (.A(net543),
    .B(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__a21oi_1 _09958_ (.A1(net543),
    .A2(_04641_),
    .B1(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__o21ai_0 _09959_ (.A1(\core.CPU_Xreg_value_a4[0][29] ),
    .A2(net470),
    .B1(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__nor2_1 _09960_ (.A(_03506_),
    .B(_03520_),
    .Y(_04646_));
 sky130_fd_sc_hd__nand2_1 _09961_ (.A(_04646_),
    .B(net432),
    .Y(_04647_));
 sky130_fd_sc_hd__o21ai_0 _09962_ (.A1(net432),
    .A2(_04645_),
    .B1(_04647_),
    .Y(\core.CPU_src1_value_a2[29] ));
 sky130_fd_sc_hd__nand3_1 _09963_ (.A(net593),
    .B(net598),
    .C(net618),
    .Y(_04648_));
 sky130_fd_sc_hd__o21ai_0 _09964_ (.A1(net543),
    .A2(\core.CPU_Xreg_value_a4[16][2] ),
    .B1(net542),
    .Y(_04649_));
 sky130_fd_sc_hd__mux4_2 _09965_ (.A0(\core.CPU_Xreg_value_a4[10][2] ),
    .A1(\core.CPU_Xreg_value_a4[11][2] ),
    .A2(\core.CPU_Xreg_value_a4[26][2] ),
    .A3(\core.CPU_Xreg_value_a4[27][2] ),
    .S0(net598),
    .S1(net593),
    .X(_04650_));
 sky130_fd_sc_hd__nor2_1 _09966_ (.A(net544),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__a31oi_1 _09967_ (.A1(net544),
    .A2(_04648_),
    .A3(_04649_),
    .B1(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__or3_1 _09968_ (.A(net596),
    .B(net593),
    .C(\core.CPU_Xreg_value_a4[0][2] ),
    .X(_04653_));
 sky130_fd_sc_hd__a21oi_1 _09969_ (.A1(\core.CPU_Xreg_value_a4[1][2] ),
    .A2(_04428_),
    .B1(_04652_),
    .Y(_04654_));
 sky130_fd_sc_hd__nor2_1 _09970_ (.A(net542),
    .B(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__a211oi_2 _09971_ (.A1(_04652_),
    .A2(_04653_),
    .B1(_04655_),
    .C1(net434),
    .Y(_04656_));
 sky130_fd_sc_hd__a21oi_1 _09972_ (.A1(_03535_),
    .A2(net432),
    .B1(net387),
    .Y(\core.CPU_src1_value_a2[2] ));
 sky130_fd_sc_hd__o21ai_0 _09973_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[1][30] ),
    .B1(net543),
    .Y(_04657_));
 sky130_fd_sc_hd__nand2_1 _09974_ (.A(net542),
    .B(\core.CPU_Xreg_value_a4[16][30] ),
    .Y(_04658_));
 sky130_fd_sc_hd__a21oi_1 _09975_ (.A1(_04657_),
    .A2(_04658_),
    .B1(net595),
    .Y(_04659_));
 sky130_fd_sc_hd__mux2_2 _09976_ (.A0(\core.CPU_Xreg_value_a4[11][30] ),
    .A1(\core.CPU_Xreg_value_a4[27][30] ),
    .S(net594),
    .X(_04660_));
 sky130_fd_sc_hd__a221oi_1 _09977_ (.A1(\core.CPU_Xreg_value_a4[17][30] ),
    .A2(net472),
    .B1(_04660_),
    .B2(net595),
    .C1(net542),
    .Y(_04661_));
 sky130_fd_sc_hd__a221oi_1 _09978_ (.A1(net543),
    .A2(\core.CPU_Xreg_value_a4[10][30] ),
    .B1(net466),
    .B2(\core.CPU_Xreg_value_a4[26][30] ),
    .C1(net597),
    .Y(_04662_));
 sky130_fd_sc_hd__nor2_1 _09979_ (.A(_04661_),
    .B(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__o22ai_1 _09980_ (.A1(\core.CPU_Xreg_value_a4[0][30] ),
    .A2(net470),
    .B1(_04659_),
    .B2(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__a21oi_1 _09981_ (.A1(net611),
    .A2(_03567_),
    .B1(_03576_),
    .Y(_04665_));
 sky130_fd_sc_hd__mux2i_1 _09982_ (.A0(_04664_),
    .A1(_04665_),
    .S(net433),
    .Y(\core.CPU_src1_value_a2[30] ));
 sky130_fd_sc_hd__a21oi_1 _09983_ (.A1(_02517_),
    .A2(net546),
    .B1(net611),
    .Y(_04666_));
 sky130_fd_sc_hd__nand4_1 _09984_ (.A(net547),
    .B(_03590_),
    .C(_03596_),
    .D(_03600_),
    .Y(_04667_));
 sky130_fd_sc_hd__nor2_1 _09985_ (.A(_01155_),
    .B(_02804_),
    .Y(_04668_));
 sky130_fd_sc_hd__nor2_1 _09986_ (.A(_03584_),
    .B(_02804_),
    .Y(_04669_));
 sky130_fd_sc_hd__inv_1 _09987_ (.A(_00200_),
    .Y(_04670_));
 sky130_fd_sc_hd__a21oi_1 _09988_ (.A1(_04670_),
    .A2(_03618_),
    .B1(_00201_),
    .Y(_04671_));
 sky130_fd_sc_hd__mux2i_1 _09989_ (.A0(_04668_),
    .A1(_04669_),
    .S(_04671_),
    .Y(_04672_));
 sky130_fd_sc_hd__o211ai_1 _09990_ (.A1(_04666_),
    .A2(_03607_),
    .B1(_04667_),
    .C1(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__mux4_2 _09991_ (.A0(\core.CPU_Xreg_value_a4[16][31] ),
    .A1(\core.CPU_Xreg_value_a4[17][31] ),
    .A2(\core.CPU_Xreg_value_a4[26][31] ),
    .A3(\core.CPU_Xreg_value_a4[27][31] ),
    .S0(net598),
    .S1(net596),
    .X(_04674_));
 sky130_fd_sc_hd__mux2i_1 _09992_ (.A0(\core.CPU_Xreg_value_a4[10][31] ),
    .A1(\core.CPU_Xreg_value_a4[11][31] ),
    .S(net598),
    .Y(_04675_));
 sky130_fd_sc_hd__nor2_1 _09993_ (.A(\core.CPU_Xreg_value_a4[1][31] ),
    .B(net465),
    .Y(_04676_));
 sky130_fd_sc_hd__a211oi_1 _09994_ (.A1(net596),
    .A2(_04675_),
    .B1(_04676_),
    .C1(\core.CPU_rf_rd_index1_a2[4] ),
    .Y(_04677_));
 sky130_fd_sc_hd__a21oi_1 _09995_ (.A1(\core.CPU_rf_rd_index1_a2[4] ),
    .A2(_04674_),
    .B1(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__nor2_1 _09996_ (.A(\core.CPU_Xreg_value_a4[0][31] ),
    .B(net470),
    .Y(_04679_));
 sky130_fd_sc_hd__nor3_1 _09997_ (.A(net433),
    .B(net401),
    .C(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__a21o_1 _09998_ (.A1(net433),
    .A2(_04673_),
    .B1(_04680_),
    .X(\core.CPU_src1_value_a2[31] ));
 sky130_fd_sc_hd__mux2_2 _09999_ (.A0(\core.CPU_Xreg_value_a4[10][3] ),
    .A1(\core.CPU_Xreg_value_a4[11][3] ),
    .S(net598),
    .X(_04681_));
 sky130_fd_sc_hd__o22ai_1 _10000_ (.A1(\core.CPU_Xreg_value_a4[1][3] ),
    .A2(net465),
    .B1(_04681_),
    .B2(net544),
    .Y(_04682_));
 sky130_fd_sc_hd__mux4_2 _10001_ (.A0(\core.CPU_Xreg_value_a4[16][3] ),
    .A1(\core.CPU_Xreg_value_a4[17][3] ),
    .A2(\core.CPU_Xreg_value_a4[26][3] ),
    .A3(\core.CPU_Xreg_value_a4[27][3] ),
    .S0(net598),
    .S1(net596),
    .X(_04683_));
 sky130_fd_sc_hd__nor2_1 _10002_ (.A(net543),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__a21oi_1 _10003_ (.A1(net543),
    .A2(_04682_),
    .B1(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__o21ai_0 _10004_ (.A1(\core.CPU_Xreg_value_a4[0][3] ),
    .A2(net469),
    .B1(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand2_1 _10005_ (.A(net372),
    .B(net434),
    .Y(_04687_));
 sky130_fd_sc_hd__o21ai_0 _10006_ (.A1(net434),
    .A2(_04686_),
    .B1(_04687_),
    .Y(\core.CPU_src1_value_a2[3] ));
 sky130_fd_sc_hd__nand3_1 _10007_ (.A(\core.CPU_rf_rd_index1_a2[4] ),
    .B(net598),
    .C(net617),
    .Y(_04688_));
 sky130_fd_sc_hd__o21ai_0 _10008_ (.A1(net543),
    .A2(\core.CPU_Xreg_value_a4[16][4] ),
    .B1(net542),
    .Y(_04689_));
 sky130_fd_sc_hd__mux4_2 _10009_ (.A0(\core.CPU_Xreg_value_a4[10][4] ),
    .A1(\core.CPU_Xreg_value_a4[11][4] ),
    .A2(\core.CPU_Xreg_value_a4[26][4] ),
    .A3(\core.CPU_Xreg_value_a4[27][4] ),
    .S0(net598),
    .S1(\core.CPU_rf_rd_index1_a2[4] ),
    .X(_04690_));
 sky130_fd_sc_hd__nor2_1 _10010_ (.A(net544),
    .B(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__a31o_2 _10011_ (.A1(net544),
    .A2(_04688_),
    .A3(_04689_),
    .B1(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__nor3_1 _10012_ (.A(net596),
    .B(net593),
    .C(\core.CPU_Xreg_value_a4[0][4] ),
    .Y(_04693_));
 sky130_fd_sc_hd__nor2_1 _10013_ (.A(_04692_),
    .B(_04693_),
    .Y(_04694_));
 sky130_fd_sc_hd__nand2_1 _10014_ (.A(\core.CPU_Xreg_value_a4[1][4] ),
    .B(_04428_),
    .Y(_04695_));
 sky130_fd_sc_hd__a21oi_1 _10015_ (.A1(_04692_),
    .A2(_04695_),
    .B1(net542),
    .Y(_04696_));
 sky130_fd_sc_hd__nor3_2 _10016_ (.A(net434),
    .B(_04694_),
    .C(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__a21oi_1 _10017_ (.A1(_03659_),
    .A2(net432),
    .B1(net400),
    .Y(\core.CPU_src1_value_a2[4] ));
 sky130_fd_sc_hd__mux2i_1 _10018_ (.A0(\core.CPU_Xreg_value_a4[26][5] ),
    .A1(\core.CPU_Xreg_value_a4[27][5] ),
    .S(net598),
    .Y(_04698_));
 sky130_fd_sc_hd__nand2_1 _10019_ (.A(\core.CPU_Xreg_value_a4[11][5] ),
    .B(net468),
    .Y(_04699_));
 sky130_fd_sc_hd__o21ai_0 _10020_ (.A1(net543),
    .A2(_04698_),
    .B1(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__o21a_1 _10021_ (.A1(net543),
    .A2(\core.CPU_Xreg_value_a4[16][5] ),
    .B1(net544),
    .X(_04701_));
 sky130_fd_sc_hd__a21oi_1 _10022_ (.A1(net543),
    .A2(\core.CPU_Xreg_value_a4[10][5] ),
    .B1(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__mux2i_1 _10023_ (.A0(\core.CPU_Xreg_value_a4[1][5] ),
    .A1(\core.CPU_Xreg_value_a4[17][5] ),
    .S(net593),
    .Y(_04703_));
 sky130_fd_sc_hd__o22ai_1 _10024_ (.A1(net598),
    .A2(_04702_),
    .B1(_04703_),
    .B2(net465),
    .Y(_04704_));
 sky130_fd_sc_hd__a21oi_1 _10025_ (.A1(net596),
    .A2(_04700_),
    .B1(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__nor2_1 _10026_ (.A(\core.CPU_Xreg_value_a4[0][5] ),
    .B(net469),
    .Y(_04706_));
 sky130_fd_sc_hd__nor2_1 _10027_ (.A(_04705_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__nor2_1 _10028_ (.A(net434),
    .B(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__a21oi_1 _10029_ (.A1(_03675_),
    .A2(net432),
    .B1(_04708_),
    .Y(\core.CPU_src1_value_a2[5] ));
 sky130_fd_sc_hd__mux2i_1 _10030_ (.A0(\core.CPU_Xreg_value_a4[26][6] ),
    .A1(\core.CPU_Xreg_value_a4[27][6] ),
    .S(\core.CPU_rf_rd_index1_a2[0] ),
    .Y(_04709_));
 sky130_fd_sc_hd__nand2_1 _10031_ (.A(\core.CPU_Xreg_value_a4[16][6] ),
    .B(_04479_),
    .Y(_04710_));
 sky130_fd_sc_hd__o21ai_0 _10032_ (.A1(net545),
    .A2(_04709_),
    .B1(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__mux2_2 _10033_ (.A0(\core.CPU_Xreg_value_a4[10][6] ),
    .A1(\core.CPU_Xreg_value_a4[11][6] ),
    .S(\core.CPU_rf_rd_index1_a2[0] ),
    .X(_04712_));
 sky130_fd_sc_hd__nand2_1 _10034_ (.A(\core.CPU_rf_rd_index1_a2[0] ),
    .B(\core.CPU_Xreg_value_a4[17][6] ),
    .Y(_04713_));
 sky130_fd_sc_hd__nor2_1 _10035_ (.A(\core.CPU_Xreg_value_a4[1][6] ),
    .B(_04451_),
    .Y(_04714_));
 sky130_fd_sc_hd__a211oi_1 _10036_ (.A1(net593),
    .A2(_04713_),
    .B1(_04714_),
    .C1(net596),
    .Y(_04715_));
 sky130_fd_sc_hd__a221o_1 _10037_ (.A1(net593),
    .A2(_04711_),
    .B1(_04712_),
    .B2(_04484_),
    .C1(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__o21ai_0 _10038_ (.A1(\core.CPU_Xreg_value_a4[0][6] ),
    .A2(net469),
    .B1(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__mux2i_1 _10039_ (.A0(net386),
    .A1(_03694_),
    .S(net432),
    .Y(\core.CPU_src1_value_a2[6] ));
 sky130_fd_sc_hd__mux2_2 _10040_ (.A0(\core.CPU_Xreg_value_a4[10][7] ),
    .A1(\core.CPU_Xreg_value_a4[11][7] ),
    .S(net597),
    .X(_04718_));
 sky130_fd_sc_hd__o22ai_1 _10041_ (.A1(\core.CPU_Xreg_value_a4[1][7] ),
    .A2(net465),
    .B1(_04718_),
    .B2(net545),
    .Y(_04719_));
 sky130_fd_sc_hd__mux4_2 _10042_ (.A0(\core.CPU_Xreg_value_a4[16][7] ),
    .A1(\core.CPU_Xreg_value_a4[17][7] ),
    .A2(\core.CPU_Xreg_value_a4[26][7] ),
    .A3(\core.CPU_Xreg_value_a4[27][7] ),
    .S0(net597),
    .S1(net595),
    .X(_04720_));
 sky130_fd_sc_hd__nor2_1 _10043_ (.A(net543),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__a21oi_1 _10044_ (.A1(net543),
    .A2(_04719_),
    .B1(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__o21ai_0 _10045_ (.A1(\core.CPU_Xreg_value_a4[0][7] ),
    .A2(net470),
    .B1(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__nand2_1 _10046_ (.A(_03706_),
    .B(net432),
    .Y(_04724_));
 sky130_fd_sc_hd__o21ai_0 _10047_ (.A1(net432),
    .A2(net399),
    .B1(_04724_),
    .Y(\core.CPU_src1_value_a2[7] ));
 sky130_fd_sc_hd__mux2_2 _10048_ (.A0(\core.CPU_Xreg_value_a4[26][8] ),
    .A1(\core.CPU_Xreg_value_a4[27][8] ),
    .S(net597),
    .X(_04725_));
 sky130_fd_sc_hd__a22oi_1 _10049_ (.A1(\core.CPU_Xreg_value_a4[11][8] ),
    .A2(net468),
    .B1(_04725_),
    .B2(net594),
    .Y(_04726_));
 sky130_fd_sc_hd__a21oi_1 _10050_ (.A1(net597),
    .A2(_04008_),
    .B1(net595),
    .Y(_04727_));
 sky130_fd_sc_hd__a21oi_1 _10051_ (.A1(net542),
    .A2(\core.CPU_Xreg_value_a4[10][8] ),
    .B1(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__mux2_2 _10052_ (.A0(\core.CPU_Xreg_value_a4[16][8] ),
    .A1(\core.CPU_Xreg_value_a4[17][8] ),
    .S(net597),
    .X(_04729_));
 sky130_fd_sc_hd__nand2_1 _10053_ (.A(net472),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__o221ai_1 _10054_ (.A1(net545),
    .A2(_04726_),
    .B1(_04728_),
    .B2(net594),
    .C1(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__o21ai_0 _10055_ (.A1(\core.CPU_Xreg_value_a4[0][8] ),
    .A2(net470),
    .B1(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__or2_2 _10056_ (.A(_03711_),
    .B(_03722_),
    .X(_04733_));
 sky130_fd_sc_hd__nand2_1 _10057_ (.A(_04733_),
    .B(net433),
    .Y(_04734_));
 sky130_fd_sc_hd__o21ai_0 _10058_ (.A1(net433),
    .A2(net398),
    .B1(_04734_),
    .Y(\core.CPU_src1_value_a2[8] ));
 sky130_fd_sc_hd__mux4_2 _10059_ (.A0(\core.CPU_Xreg_value_a4[10][9] ),
    .A1(\core.CPU_Xreg_value_a4[11][9] ),
    .A2(\core.CPU_Xreg_value_a4[26][9] ),
    .A3(\core.CPU_Xreg_value_a4[27][9] ),
    .S0(net597),
    .S1(net594),
    .X(_04735_));
 sky130_fd_sc_hd__mux4_2 _10060_ (.A0(\core.CPU_Xreg_value_a4[0][9] ),
    .A1(\core.CPU_Xreg_value_a4[1][9] ),
    .A2(\core.CPU_Xreg_value_a4[16][9] ),
    .A3(\core.CPU_Xreg_value_a4[17][9] ),
    .S0(net597),
    .S1(net594),
    .X(_04736_));
 sky130_fd_sc_hd__mux2i_1 _10061_ (.A0(_04735_),
    .A1(_04736_),
    .S(net545),
    .Y(_04737_));
 sky130_fd_sc_hd__nand2_1 _10062_ (.A(_03741_),
    .B(net433),
    .Y(_04738_));
 sky130_fd_sc_hd__o21ai_0 _10063_ (.A1(net433),
    .A2(net463),
    .B1(_04738_),
    .Y(\core.CPU_src1_value_a2[9] ));
 sky130_fd_sc_hd__xor2_1 _10064_ (.A(\core.CPU_rd_a3[1] ),
    .B(net590),
    .X(_04739_));
 sky130_fd_sc_hd__xor2_1 _10065_ (.A(\core.CPU_rd_a3[3] ),
    .B(net587),
    .X(_04740_));
 sky130_fd_sc_hd__xor2_1 _10068_ (.A(\core.CPU_rd_a3[0] ),
    .B(\core.CPU_rf_rd_index2_a2[0] ),
    .X(_04743_));
 sky130_fd_sc_hd__nor4_1 _10069_ (.A(\core.CPU_rd_a3[4] ),
    .B(_04739_),
    .C(_04740_),
    .D(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__nand2_2 _10070_ (.A(_02556_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__or3_1 _10073_ (.A(\core.CPU_rf_rd_index2_a2[3] ),
    .B(net591),
    .C(net589),
    .X(_04748_));
 sky130_fd_sc_hd__inv_1 _10076_ (.A(\core.CPU_rf_rd_index2_a2[1] ),
    .Y(_04751_));
 sky130_fd_sc_hd__nor2_1 _10077_ (.A(\core.CPU_rf_rd_index2_a2[3] ),
    .B(net539),
    .Y(_04752_));
 sky130_fd_sc_hd__mux2_2 _10080_ (.A0(\core.CPU_Xreg_value_a4[2][0] ),
    .A1(\core.CPU_Xreg_value_a4[3][0] ),
    .S(net592),
    .X(_04755_));
 sky130_fd_sc_hd__mux2i_1 _10083_ (.A0(\core.CPU_Xreg_value_a4[10][0] ),
    .A1(\core.CPU_Xreg_value_a4[11][0] ),
    .S(net592),
    .Y(_04758_));
 sky130_fd_sc_hd__clkinv_1 _10084_ (.A(\core.CPU_rf_rd_index2_a2[0] ),
    .Y(_04759_));
 sky130_fd_sc_hd__nor2_2 _10085_ (.A(net538),
    .B(net590),
    .Y(_04760_));
 sky130_fd_sc_hd__nand2_1 _10087_ (.A(\core.CPU_Xreg_value_a4[9][0] ),
    .B(net461),
    .Y(_04762_));
 sky130_fd_sc_hd__o21ai_0 _10088_ (.A1(net539),
    .A2(_04758_),
    .B1(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__a21oi_1 _10096_ (.A1(_04422_),
    .A2(net592),
    .B1(net587),
    .Y(_04771_));
 sky130_fd_sc_hd__a21oi_1 _10097_ (.A1(\core.CPU_Xreg_value_a4[8][0] ),
    .A2(net538),
    .B1(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__nor2_1 _10098_ (.A(net590),
    .B(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__a221o_1 _10099_ (.A1(net462),
    .A2(_04755_),
    .B1(_04763_),
    .B2(net587),
    .C1(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__o211ai_1 _10101_ (.A1(\core.CPU_Xreg_value_a4[0][0] ),
    .A2(net540),
    .B1(_04774_),
    .C1(net430),
    .Y(_04776_));
 sky130_fd_sc_hd__o21ai_1 _10102_ (.A1(net394),
    .A2(net430),
    .B1(_04776_),
    .Y(\core.CPU_src2_value_a2[0] ));
 sky130_fd_sc_hd__mux4_2 _10105_ (.A0(\core.CPU_Xreg_value_a4[0][10] ),
    .A1(\core.CPU_Xreg_value_a4[1][10] ),
    .A2(\core.CPU_Xreg_value_a4[2][10] ),
    .A3(\core.CPU_Xreg_value_a4[3][10] ),
    .S0(net592),
    .S1(net590),
    .X(_04779_));
 sky130_fd_sc_hd__mux4_2 _10108_ (.A0(\core.CPU_Xreg_value_a4[8][10] ),
    .A1(\core.CPU_Xreg_value_a4[9][10] ),
    .A2(\core.CPU_Xreg_value_a4[10][10] ),
    .A3(\core.CPU_Xreg_value_a4[11][10] ),
    .S0(net592),
    .S1(net590),
    .X(_04782_));
 sky130_fd_sc_hd__mux2_2 _10109_ (.A0(_04779_),
    .A1(_04782_),
    .S(net587),
    .X(_04783_));
 sky130_fd_sc_hd__nand2_1 _10110_ (.A(net430),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__o21ai_0 _10111_ (.A1(_02640_),
    .A2(net431),
    .B1(_04784_),
    .Y(\core.CPU_src2_value_a2[10] ));
 sky130_fd_sc_hd__mux4_2 _10113_ (.A0(\core.CPU_Xreg_value_a4[0][11] ),
    .A1(\core.CPU_Xreg_value_a4[1][11] ),
    .A2(\core.CPU_Xreg_value_a4[2][11] ),
    .A3(\core.CPU_Xreg_value_a4[3][11] ),
    .S0(net592),
    .S1(net590),
    .X(_04786_));
 sky130_fd_sc_hd__mux4_2 _10115_ (.A0(\core.CPU_Xreg_value_a4[8][11] ),
    .A1(\core.CPU_Xreg_value_a4[9][11] ),
    .A2(\core.CPU_Xreg_value_a4[10][11] ),
    .A3(\core.CPU_Xreg_value_a4[11][11] ),
    .S0(net592),
    .S1(net590),
    .X(_04788_));
 sky130_fd_sc_hd__mux2i_2 _10118_ (.A0(_04786_),
    .A1(_04788_),
    .S(net587),
    .Y(_04791_));
 sky130_fd_sc_hd__nor2_1 _10120_ (.A(_02717_),
    .B(net431),
    .Y(_04793_));
 sky130_fd_sc_hd__a21oi_1 _10121_ (.A1(net431),
    .A2(net460),
    .B1(_04793_),
    .Y(\core.CPU_src2_value_a2[11] ));
 sky130_fd_sc_hd__mux4_2 _10122_ (.A0(\core.CPU_Xreg_value_a4[0][12] ),
    .A1(\core.CPU_Xreg_value_a4[1][12] ),
    .A2(\core.CPU_Xreg_value_a4[2][12] ),
    .A3(\core.CPU_Xreg_value_a4[3][12] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(net589),
    .X(_04794_));
 sky130_fd_sc_hd__nor2_1 _10125_ (.A(net588),
    .B(_04794_),
    .Y(_04797_));
 sky130_fd_sc_hd__mux2_2 _10127_ (.A0(\core.CPU_Xreg_value_a4[10][12] ),
    .A1(\core.CPU_Xreg_value_a4[11][12] ),
    .S(\core.CPU_rf_rd_index2_a2[0] ),
    .X(_04799_));
 sky130_fd_sc_hd__nand2_1 _10128_ (.A(\core.CPU_Xreg_value_a4[9][12] ),
    .B(net461),
    .Y(_04800_));
 sky130_fd_sc_hd__nand2_1 _10129_ (.A(net588),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__a21oi_1 _10130_ (.A1(net589),
    .A2(_04799_),
    .B1(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__nor2_1 _10132_ (.A(\core.CPU_rf_rd_index2_a2[0] ),
    .B(net589),
    .Y(_04804_));
 sky130_fd_sc_hd__nand2_1 _10133_ (.A(\core.CPU_Xreg_value_a4[8][12] ),
    .B(net537),
    .Y(_04805_));
 sky130_fd_sc_hd__o21ai_0 _10134_ (.A1(_04797_),
    .A2(_04802_),
    .B1(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__o311ai_1 _10136_ (.A1(\core.CPU_Xreg_value_a4[0][12] ),
    .A2(net588),
    .A3(_04794_),
    .B1(_04806_),
    .C1(net430),
    .Y(_04808_));
 sky130_fd_sc_hd__o21ai_0 _10137_ (.A1(_04476_),
    .A2(net431),
    .B1(net379),
    .Y(\core.CPU_src2_value_a2[12] ));
 sky130_fd_sc_hd__nor2b_1 _10139_ (.A(net589),
    .B_N(net588),
    .Y(_04810_));
 sky130_fd_sc_hd__a22oi_1 _10140_ (.A1(\core.CPU_Xreg_value_a4[2][13] ),
    .A2(net462),
    .B1(_04810_),
    .B2(\core.CPU_Xreg_value_a4[8][13] ),
    .Y(_04811_));
 sky130_fd_sc_hd__nor2_1 _10141_ (.A(\core.CPU_rf_rd_index2_a2[3] ),
    .B(net589),
    .Y(_04812_));
 sky130_fd_sc_hd__o21ai_0 _10142_ (.A1(\core.CPU_Xreg_value_a4[1][13] ),
    .A2(net538),
    .B1(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__mux2_2 _10143_ (.A0(\core.CPU_Xreg_value_a4[3][13] ),
    .A1(\core.CPU_Xreg_value_a4[11][13] ),
    .S(\core.CPU_rf_rd_index2_a2[3] ),
    .X(_04814_));
 sky130_fd_sc_hd__nand3_1 _10144_ (.A(net591),
    .B(net589),
    .C(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nor2_1 _10145_ (.A(net591),
    .B(net539),
    .Y(_04816_));
 sky130_fd_sc_hd__a22o_1 _10146_ (.A1(\core.CPU_Xreg_value_a4[9][13] ),
    .A2(net461),
    .B1(_04816_),
    .B2(\core.CPU_Xreg_value_a4[10][13] ),
    .X(_04817_));
 sky130_fd_sc_hd__nand2_1 _10147_ (.A(\core.CPU_rf_rd_index2_a2[3] ),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__o2111ai_1 _10148_ (.A1(net591),
    .A2(_04811_),
    .B1(_04813_),
    .C1(_04815_),
    .D1(_04818_),
    .Y(_04819_));
 sky130_fd_sc_hd__o211ai_1 _10149_ (.A1(\core.CPU_Xreg_value_a4[0][13] ),
    .A2(net540),
    .B1(_04819_),
    .C1(net430),
    .Y(_04820_));
 sky130_fd_sc_hd__o21ai_0 _10150_ (.A1(_02810_),
    .A2(net430),
    .B1(_04820_),
    .Y(\core.CPU_src2_value_a2[13] ));
 sky130_fd_sc_hd__mux4_2 _10151_ (.A0(\core.CPU_Xreg_value_a4[0][14] ),
    .A1(\core.CPU_Xreg_value_a4[1][14] ),
    .A2(\core.CPU_Xreg_value_a4[2][14] ),
    .A3(\core.CPU_Xreg_value_a4[3][14] ),
    .S0(net592),
    .S1(net590),
    .X(_04821_));
 sky130_fd_sc_hd__mux4_2 _10152_ (.A0(\core.CPU_Xreg_value_a4[8][14] ),
    .A1(\core.CPU_Xreg_value_a4[9][14] ),
    .A2(\core.CPU_Xreg_value_a4[10][14] ),
    .A3(\core.CPU_Xreg_value_a4[11][14] ),
    .S0(net592),
    .S1(net590),
    .X(_04822_));
 sky130_fd_sc_hd__mux2_2 _10153_ (.A0(_04821_),
    .A1(_04822_),
    .S(net587),
    .X(_04823_));
 sky130_fd_sc_hd__nand2_1 _10154_ (.A(net430),
    .B(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__o21ai_0 _10155_ (.A1(_02866_),
    .A2(net431),
    .B1(_04824_),
    .Y(\core.CPU_src2_value_a2[14] ));
 sky130_fd_sc_hd__mux2_2 _10156_ (.A0(\core.CPU_Xreg_value_a4[9][15] ),
    .A1(\core.CPU_Xreg_value_a4[11][15] ),
    .S(net589),
    .X(_04825_));
 sky130_fd_sc_hd__a22oi_1 _10157_ (.A1(\core.CPU_Xreg_value_a4[3][15] ),
    .A2(_04752_),
    .B1(_04825_),
    .B2(net588),
    .Y(_04826_));
 sky130_fd_sc_hd__o21ai_0 _10159_ (.A1(\core.CPU_Xreg_value_a4[2][15] ),
    .A2(net539),
    .B1(net538),
    .Y(_04828_));
 sky130_fd_sc_hd__a21boi_0 _10160_ (.A1(\core.CPU_Xreg_value_a4[1][15] ),
    .A2(net539),
    .B1_N(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__mux2i_1 _10161_ (.A0(\core.CPU_Xreg_value_a4[8][15] ),
    .A1(\core.CPU_Xreg_value_a4[10][15] ),
    .S(net589),
    .Y(_04830_));
 sky130_fd_sc_hd__nand2_1 _10162_ (.A(net587),
    .B(net538),
    .Y(_04831_));
 sky130_fd_sc_hd__o22a_1 _10163_ (.A1(\core.CPU_rf_rd_index2_a2[3] ),
    .A2(_04829_),
    .B1(_04830_),
    .B2(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__o21ai_0 _10164_ (.A1(net538),
    .A2(_04826_),
    .B1(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__o211ai_1 _10165_ (.A1(\core.CPU_Xreg_value_a4[0][15] ),
    .A2(net540),
    .B1(_04833_),
    .C1(net430),
    .Y(_04834_));
 sky130_fd_sc_hd__o21ai_0 _10166_ (.A1(_02909_),
    .A2(net430),
    .B1(_04834_),
    .Y(\core.CPU_src2_value_a2[15] ));
 sky130_fd_sc_hd__mux4_2 _10167_ (.A0(\core.CPU_Xreg_value_a4[0][16] ),
    .A1(\core.CPU_Xreg_value_a4[1][16] ),
    .A2(\core.CPU_Xreg_value_a4[2][16] ),
    .A3(\core.CPU_Xreg_value_a4[3][16] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(net589),
    .X(_04835_));
 sky130_fd_sc_hd__or3_1 _10168_ (.A(\core.CPU_Xreg_value_a4[0][16] ),
    .B(net588),
    .C(_04835_),
    .X(_04836_));
 sky130_fd_sc_hd__mux2_2 _10169_ (.A0(\core.CPU_Xreg_value_a4[10][16] ),
    .A1(\core.CPU_Xreg_value_a4[11][16] ),
    .S(\core.CPU_rf_rd_index2_a2[0] ),
    .X(_04837_));
 sky130_fd_sc_hd__nand2_1 _10170_ (.A(net589),
    .B(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__nand2_1 _10171_ (.A(\core.CPU_Xreg_value_a4[9][16] ),
    .B(net461),
    .Y(_04839_));
 sky130_fd_sc_hd__nor2_1 _10172_ (.A(net588),
    .B(_04835_),
    .Y(_04840_));
 sky130_fd_sc_hd__a31oi_1 _10173_ (.A1(net588),
    .A2(_04838_),
    .A3(_04839_),
    .B1(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__a31oi_1 _10174_ (.A1(\core.CPU_Xreg_value_a4[8][16] ),
    .A2(net537),
    .A3(_04836_),
    .B1(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__nor2_1 _10175_ (.A(_02956_),
    .B(net430),
    .Y(_04843_));
 sky130_fd_sc_hd__a21oi_1 _10176_ (.A1(net430),
    .A2(_04842_),
    .B1(_04843_),
    .Y(\core.CPU_src2_value_a2[16] ));
 sky130_fd_sc_hd__mux2_2 _10177_ (.A0(\core.CPU_Xreg_value_a4[9][17] ),
    .A1(\core.CPU_Xreg_value_a4[11][17] ),
    .S(net589),
    .X(_04844_));
 sky130_fd_sc_hd__a22o_1 _10178_ (.A1(\core.CPU_Xreg_value_a4[3][17] ),
    .A2(net462),
    .B1(_04844_),
    .B2(net588),
    .X(_04845_));
 sky130_fd_sc_hd__inv_1 _10179_ (.A(\core.CPU_Xreg_value_a4[2][17] ),
    .Y(_04846_));
 sky130_fd_sc_hd__mux2i_1 _10180_ (.A0(\core.CPU_Xreg_value_a4[8][17] ),
    .A1(\core.CPU_Xreg_value_a4[10][17] ),
    .S(net589),
    .Y(_04847_));
 sky130_fd_sc_hd__a221oi_1 _10181_ (.A1(_04846_),
    .A2(net462),
    .B1(_04847_),
    .B2(net588),
    .C1(net591),
    .Y(_04848_));
 sky130_fd_sc_hd__a221o_1 _10182_ (.A1(\core.CPU_Xreg_value_a4[1][17] ),
    .A2(_04812_),
    .B1(_04845_),
    .B2(net591),
    .C1(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__o211ai_1 _10183_ (.A1(\core.CPU_Xreg_value_a4[0][17] ),
    .A2(net540),
    .B1(_04849_),
    .C1(net430),
    .Y(_04850_));
 sky130_fd_sc_hd__o21ai_0 _10184_ (.A1(_03003_),
    .A2(net430),
    .B1(_04850_),
    .Y(\core.CPU_src2_value_a2[17] ));
 sky130_fd_sc_hd__mux4_2 _10185_ (.A0(\core.CPU_Xreg_value_a4[0][18] ),
    .A1(\core.CPU_Xreg_value_a4[1][18] ),
    .A2(\core.CPU_Xreg_value_a4[2][18] ),
    .A3(\core.CPU_Xreg_value_a4[3][18] ),
    .S0(net591),
    .S1(net589),
    .X(_04851_));
 sky130_fd_sc_hd__mux4_2 _10186_ (.A0(\core.CPU_Xreg_value_a4[8][18] ),
    .A1(\core.CPU_Xreg_value_a4[9][18] ),
    .A2(\core.CPU_Xreg_value_a4[10][18] ),
    .A3(\core.CPU_Xreg_value_a4[11][18] ),
    .S0(net591),
    .S1(net589),
    .X(_04852_));
 sky130_fd_sc_hd__mux2_2 _10187_ (.A0(_04851_),
    .A1(_04852_),
    .S(net588),
    .X(_04853_));
 sky130_fd_sc_hd__nand2_1 _10188_ (.A(net430),
    .B(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__o21ai_0 _10189_ (.A1(net359),
    .A2(net430),
    .B1(_04854_),
    .Y(\core.CPU_src2_value_a2[18] ));
 sky130_fd_sc_hd__mux4_2 _10190_ (.A0(\core.CPU_Xreg_value_a4[0][19] ),
    .A1(\core.CPU_Xreg_value_a4[1][19] ),
    .A2(\core.CPU_Xreg_value_a4[2][19] ),
    .A3(\core.CPU_Xreg_value_a4[3][19] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(\core.CPU_rf_rd_index2_a2[1] ),
    .X(_04855_));
 sky130_fd_sc_hd__nor2_1 _10191_ (.A(net588),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__mux2_2 _10192_ (.A0(\core.CPU_Xreg_value_a4[10][19] ),
    .A1(\core.CPU_Xreg_value_a4[11][19] ),
    .S(\core.CPU_rf_rd_index2_a2[0] ),
    .X(_04857_));
 sky130_fd_sc_hd__nand2_1 _10193_ (.A(\core.CPU_Xreg_value_a4[9][19] ),
    .B(net461),
    .Y(_04858_));
 sky130_fd_sc_hd__nand2_1 _10194_ (.A(net588),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__a21oi_1 _10195_ (.A1(\core.CPU_rf_rd_index2_a2[1] ),
    .A2(_04857_),
    .B1(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__nand2_1 _10196_ (.A(\core.CPU_Xreg_value_a4[8][19] ),
    .B(net537),
    .Y(_04861_));
 sky130_fd_sc_hd__o21ai_0 _10197_ (.A1(_04856_),
    .A2(_04860_),
    .B1(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__o311ai_0 _10198_ (.A1(\core.CPU_Xreg_value_a4[0][19] ),
    .A2(net588),
    .A3(_04855_),
    .B1(_04862_),
    .C1(net430),
    .Y(_04863_));
 sky130_fd_sc_hd__o21ai_0 _10199_ (.A1(_04534_),
    .A2(net431),
    .B1(net378),
    .Y(\core.CPU_src2_value_a2[19] ));
 sky130_fd_sc_hd__mux4_2 _10200_ (.A0(\core.CPU_Xreg_value_a4[0][1] ),
    .A1(\core.CPU_Xreg_value_a4[1][1] ),
    .A2(\core.CPU_Xreg_value_a4[2][1] ),
    .A3(\core.CPU_Xreg_value_a4[3][1] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(\core.CPU_rf_rd_index2_a2[1] ),
    .X(_04864_));
 sky130_fd_sc_hd__or3_1 _10201_ (.A(\core.CPU_Xreg_value_a4[0][1] ),
    .B(net587),
    .C(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__mux2_2 _10202_ (.A0(\core.CPU_Xreg_value_a4[10][1] ),
    .A1(\core.CPU_Xreg_value_a4[11][1] ),
    .S(\core.CPU_rf_rd_index2_a2[0] ),
    .X(_04866_));
 sky130_fd_sc_hd__nand2_1 _10203_ (.A(\core.CPU_rf_rd_index2_a2[1] ),
    .B(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__nand2_1 _10204_ (.A(\core.CPU_Xreg_value_a4[9][1] ),
    .B(net461),
    .Y(_04868_));
 sky130_fd_sc_hd__nor2_1 _10205_ (.A(net587),
    .B(_04864_),
    .Y(_04869_));
 sky130_fd_sc_hd__a31oi_1 _10206_ (.A1(net587),
    .A2(_04867_),
    .A3(_04868_),
    .B1(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__a31oi_1 _10207_ (.A1(\core.CPU_Xreg_value_a4[8][1] ),
    .A2(net537),
    .A3(_04865_),
    .B1(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__nor2_1 _10208_ (.A(_03099_),
    .B(net431),
    .Y(_04872_));
 sky130_fd_sc_hd__a21oi_1 _10209_ (.A1(net431),
    .A2(net397),
    .B1(_04872_),
    .Y(\core.CPU_src2_value_a2[1] ));
 sky130_fd_sc_hd__mux4_2 _10210_ (.A0(\core.CPU_Xreg_value_a4[0][20] ),
    .A1(\core.CPU_Xreg_value_a4[1][20] ),
    .A2(\core.CPU_Xreg_value_a4[2][20] ),
    .A3(\core.CPU_Xreg_value_a4[3][20] ),
    .S0(net592),
    .S1(net590),
    .X(_04873_));
 sky130_fd_sc_hd__or3_1 _10211_ (.A(\core.CPU_Xreg_value_a4[0][20] ),
    .B(net587),
    .C(_04873_),
    .X(_04874_));
 sky130_fd_sc_hd__mux2_2 _10212_ (.A0(\core.CPU_Xreg_value_a4[10][20] ),
    .A1(\core.CPU_Xreg_value_a4[11][20] ),
    .S(net592),
    .X(_04875_));
 sky130_fd_sc_hd__nand2_1 _10213_ (.A(net590),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__nand2_1 _10214_ (.A(\core.CPU_Xreg_value_a4[9][20] ),
    .B(_04760_),
    .Y(_04877_));
 sky130_fd_sc_hd__nor2_1 _10215_ (.A(net587),
    .B(_04873_),
    .Y(_04878_));
 sky130_fd_sc_hd__a31oi_1 _10216_ (.A1(net587),
    .A2(_04876_),
    .A3(_04877_),
    .B1(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__a31oi_2 _10217_ (.A1(\core.CPU_Xreg_value_a4[8][20] ),
    .A2(net537),
    .A3(_04874_),
    .B1(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__nor2_1 _10218_ (.A(_03141_),
    .B(net431),
    .Y(_04881_));
 sky130_fd_sc_hd__a21oi_1 _10219_ (.A1(net431),
    .A2(net396),
    .B1(_04881_),
    .Y(\core.CPU_src2_value_a2[20] ));
 sky130_fd_sc_hd__mux4_2 _10220_ (.A0(\core.CPU_Xreg_value_a4[0][21] ),
    .A1(\core.CPU_Xreg_value_a4[1][21] ),
    .A2(\core.CPU_Xreg_value_a4[2][21] ),
    .A3(\core.CPU_Xreg_value_a4[3][21] ),
    .S0(net592),
    .S1(net590),
    .X(_04882_));
 sky130_fd_sc_hd__mux4_2 _10221_ (.A0(\core.CPU_Xreg_value_a4[8][21] ),
    .A1(\core.CPU_Xreg_value_a4[9][21] ),
    .A2(\core.CPU_Xreg_value_a4[10][21] ),
    .A3(\core.CPU_Xreg_value_a4[11][21] ),
    .S0(net592),
    .S1(net590),
    .X(_04883_));
 sky130_fd_sc_hd__mux2i_2 _10222_ (.A0(_04882_),
    .A1(_04883_),
    .S(net587),
    .Y(_04884_));
 sky130_fd_sc_hd__nor2_1 _10223_ (.A(_03188_),
    .B(net431),
    .Y(_04885_));
 sky130_fd_sc_hd__a21oi_1 _10224_ (.A1(net431),
    .A2(net458),
    .B1(_04885_),
    .Y(\core.CPU_src2_value_a2[21] ));
 sky130_fd_sc_hd__mux2_2 _10225_ (.A0(\core.CPU_Xreg_value_a4[9][22] ),
    .A1(\core.CPU_Xreg_value_a4[11][22] ),
    .S(net589),
    .X(_04886_));
 sky130_fd_sc_hd__a22oi_1 _10226_ (.A1(\core.CPU_Xreg_value_a4[3][22] ),
    .A2(_04752_),
    .B1(_04886_),
    .B2(net588),
    .Y(_04887_));
 sky130_fd_sc_hd__o21ai_0 _10227_ (.A1(\core.CPU_Xreg_value_a4[2][22] ),
    .A2(net539),
    .B1(net538),
    .Y(_04888_));
 sky130_fd_sc_hd__a21boi_0 _10228_ (.A1(\core.CPU_Xreg_value_a4[1][22] ),
    .A2(net539),
    .B1_N(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__mux2i_1 _10229_ (.A0(\core.CPU_Xreg_value_a4[8][22] ),
    .A1(\core.CPU_Xreg_value_a4[10][22] ),
    .S(net589),
    .Y(_04890_));
 sky130_fd_sc_hd__o22a_1 _10230_ (.A1(net588),
    .A2(_04889_),
    .B1(_04890_),
    .B2(_04831_),
    .X(_04891_));
 sky130_fd_sc_hd__o21ai_0 _10231_ (.A1(net538),
    .A2(_04887_),
    .B1(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__o211ai_1 _10232_ (.A1(\core.CPU_Xreg_value_a4[0][22] ),
    .A2(net540),
    .B1(_04892_),
    .C1(net430),
    .Y(_04893_));
 sky130_fd_sc_hd__o21ai_0 _10233_ (.A1(_04578_),
    .A2(net430),
    .B1(_04893_),
    .Y(\core.CPU_src2_value_a2[22] ));
 sky130_fd_sc_hd__mux2_2 _10234_ (.A0(\core.CPU_Xreg_value_a4[9][23] ),
    .A1(\core.CPU_Xreg_value_a4[11][23] ),
    .S(net589),
    .X(_04894_));
 sky130_fd_sc_hd__a22o_1 _10235_ (.A1(\core.CPU_Xreg_value_a4[3][23] ),
    .A2(net462),
    .B1(_04894_),
    .B2(\core.CPU_rf_rd_index2_a2[3] ),
    .X(_04895_));
 sky130_fd_sc_hd__inv_1 _10236_ (.A(\core.CPU_Xreg_value_a4[2][23] ),
    .Y(_04896_));
 sky130_fd_sc_hd__mux2i_1 _10237_ (.A0(\core.CPU_Xreg_value_a4[8][23] ),
    .A1(\core.CPU_Xreg_value_a4[10][23] ),
    .S(net589),
    .Y(_04897_));
 sky130_fd_sc_hd__a221oi_1 _10238_ (.A1(_04896_),
    .A2(net462),
    .B1(_04897_),
    .B2(\core.CPU_rf_rd_index2_a2[3] ),
    .C1(net591),
    .Y(_04898_));
 sky130_fd_sc_hd__a221o_1 _10239_ (.A1(\core.CPU_Xreg_value_a4[1][23] ),
    .A2(_04812_),
    .B1(_04895_),
    .B2(net591),
    .C1(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__o211ai_1 _10240_ (.A1(\core.CPU_Xreg_value_a4[0][23] ),
    .A2(net540),
    .B1(_04899_),
    .C1(net430),
    .Y(_04900_));
 sky130_fd_sc_hd__o21ai_0 _10241_ (.A1(_04579_),
    .A2(net430),
    .B1(_04900_),
    .Y(\core.CPU_src2_value_a2[23] ));
 sky130_fd_sc_hd__mux2_2 _10242_ (.A0(\core.CPU_Xreg_value_a4[9][24] ),
    .A1(\core.CPU_Xreg_value_a4[11][24] ),
    .S(net589),
    .X(_04901_));
 sky130_fd_sc_hd__a22o_1 _10243_ (.A1(\core.CPU_Xreg_value_a4[3][24] ),
    .A2(net462),
    .B1(_04901_),
    .B2(\core.CPU_rf_rd_index2_a2[3] ),
    .X(_04902_));
 sky130_fd_sc_hd__o21ai_0 _10244_ (.A1(\core.CPU_Xreg_value_a4[2][24] ),
    .A2(net539),
    .B1(net538),
    .Y(_04903_));
 sky130_fd_sc_hd__a21boi_0 _10245_ (.A1(\core.CPU_Xreg_value_a4[1][24] ),
    .A2(net539),
    .B1_N(_04903_),
    .Y(_04904_));
 sky130_fd_sc_hd__mux2i_1 _10246_ (.A0(\core.CPU_Xreg_value_a4[8][24] ),
    .A1(\core.CPU_Xreg_value_a4[10][24] ),
    .S(net589),
    .Y(_04905_));
 sky130_fd_sc_hd__o22ai_1 _10247_ (.A1(net588),
    .A2(_04904_),
    .B1(_04905_),
    .B2(_04831_),
    .Y(_04906_));
 sky130_fd_sc_hd__a21oi_1 _10248_ (.A1(net591),
    .A2(_04902_),
    .B1(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__nor2_1 _10249_ (.A(\core.CPU_Xreg_value_a4[0][24] ),
    .B(net540),
    .Y(_04908_));
 sky130_fd_sc_hd__o21ai_0 _10250_ (.A1(_04907_),
    .A2(_04908_),
    .B1(net430),
    .Y(_04909_));
 sky130_fd_sc_hd__o21a_1 _10251_ (.A1(_04589_),
    .A2(net430),
    .B1(_04909_),
    .X(\core.CPU_src2_value_a2[24] ));
 sky130_fd_sc_hd__mux4_2 _10252_ (.A0(\core.CPU_Xreg_value_a4[0][25] ),
    .A1(\core.CPU_Xreg_value_a4[1][25] ),
    .A2(\core.CPU_Xreg_value_a4[2][25] ),
    .A3(\core.CPU_Xreg_value_a4[3][25] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(\core.CPU_rf_rd_index2_a2[1] ),
    .X(_04910_));
 sky130_fd_sc_hd__mux4_2 _10253_ (.A0(\core.CPU_Xreg_value_a4[8][25] ),
    .A1(\core.CPU_Xreg_value_a4[9][25] ),
    .A2(\core.CPU_Xreg_value_a4[10][25] ),
    .A3(\core.CPU_Xreg_value_a4[11][25] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(\core.CPU_rf_rd_index2_a2[1] ),
    .X(_04911_));
 sky130_fd_sc_hd__mux2i_1 _10254_ (.A0(_04910_),
    .A1(_04911_),
    .S(net588),
    .Y(_04912_));
 sky130_fd_sc_hd__nor2_1 _10255_ (.A(_03352_),
    .B(net430),
    .Y(_04913_));
 sky130_fd_sc_hd__a21oi_1 _10256_ (.A1(net430),
    .A2(_04912_),
    .B1(_04913_),
    .Y(\core.CPU_src2_value_a2[25] ));
 sky130_fd_sc_hd__a22oi_1 _10257_ (.A1(\core.CPU_Xreg_value_a4[2][26] ),
    .A2(net462),
    .B1(_04810_),
    .B2(\core.CPU_Xreg_value_a4[8][26] ),
    .Y(_04914_));
 sky130_fd_sc_hd__nor2_1 _10258_ (.A(net591),
    .B(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__nand3b_1 _10259_ (.A_N(net588),
    .B(net591),
    .C(\core.CPU_Xreg_value_a4[3][26] ),
    .Y(_04916_));
 sky130_fd_sc_hd__mux2_2 _10260_ (.A0(\core.CPU_Xreg_value_a4[10][26] ),
    .A1(\core.CPU_Xreg_value_a4[11][26] ),
    .S(net591),
    .X(_04917_));
 sky130_fd_sc_hd__nand2_1 _10261_ (.A(net588),
    .B(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__a21oi_1 _10262_ (.A1(_04610_),
    .A2(net591),
    .B1(net588),
    .Y(_04919_));
 sky130_fd_sc_hd__a311oi_1 _10263_ (.A1(\core.CPU_Xreg_value_a4[9][26] ),
    .A2(net588),
    .A3(net591),
    .B1(net589),
    .C1(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__a31oi_1 _10264_ (.A1(net589),
    .A2(_04916_),
    .A3(_04918_),
    .B1(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__o221ai_1 _10265_ (.A1(\core.CPU_Xreg_value_a4[0][26] ),
    .A2(net540),
    .B1(_04915_),
    .B2(_04921_),
    .C1(net430),
    .Y(_04922_));
 sky130_fd_sc_hd__o21ai_0 _10266_ (.A1(_03387_),
    .A2(net430),
    .B1(_04922_),
    .Y(\core.CPU_src2_value_a2[26] ));
 sky130_fd_sc_hd__mux4_2 _10267_ (.A0(\core.CPU_Xreg_value_a4[0][27] ),
    .A1(\core.CPU_Xreg_value_a4[1][27] ),
    .A2(\core.CPU_Xreg_value_a4[2][27] ),
    .A3(\core.CPU_Xreg_value_a4[3][27] ),
    .S0(net591),
    .S1(net589),
    .X(_04923_));
 sky130_fd_sc_hd__mux4_2 _10268_ (.A0(\core.CPU_Xreg_value_a4[8][27] ),
    .A1(\core.CPU_Xreg_value_a4[9][27] ),
    .A2(\core.CPU_Xreg_value_a4[10][27] ),
    .A3(\core.CPU_Xreg_value_a4[11][27] ),
    .S0(net591),
    .S1(net589),
    .X(_04924_));
 sky130_fd_sc_hd__mux2i_1 _10269_ (.A0(_04923_),
    .A1(_04924_),
    .S(net588),
    .Y(_04925_));
 sky130_fd_sc_hd__a21oi_1 _10270_ (.A1(net367),
    .A2(_03430_),
    .B1(net430),
    .Y(_04926_));
 sky130_fd_sc_hd__a22oi_1 _10271_ (.A1(net430),
    .A2(_04925_),
    .B1(_04926_),
    .B2(net353),
    .Y(\core.CPU_src2_value_a2[27] ));
 sky130_fd_sc_hd__a22oi_1 _10272_ (.A1(\core.CPU_Xreg_value_a4[3][28] ),
    .A2(net462),
    .B1(_04810_),
    .B2(\core.CPU_Xreg_value_a4[9][28] ),
    .Y(_04927_));
 sky130_fd_sc_hd__nor2_1 _10273_ (.A(net538),
    .B(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _10274_ (.A(\core.CPU_Xreg_value_a4[11][28] ),
    .B(net591),
    .Y(_04929_));
 sky130_fd_sc_hd__o21ai_0 _10275_ (.A1(_04631_),
    .A2(net591),
    .B1(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__nor2_1 _10276_ (.A(net588),
    .B(net591),
    .Y(_04931_));
 sky130_fd_sc_hd__a22oi_1 _10277_ (.A1(net588),
    .A2(_04930_),
    .B1(_04931_),
    .B2(\core.CPU_Xreg_value_a4[2][28] ),
    .Y(_04932_));
 sky130_fd_sc_hd__nor2_1 _10278_ (.A(net539),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__inv_1 _10279_ (.A(\core.CPU_Xreg_value_a4[1][28] ),
    .Y(_04934_));
 sky130_fd_sc_hd__a21oi_1 _10280_ (.A1(_04934_),
    .A2(net591),
    .B1(net588),
    .Y(_04935_));
 sky130_fd_sc_hd__a21oi_1 _10281_ (.A1(\core.CPU_Xreg_value_a4[8][28] ),
    .A2(net538),
    .B1(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__nor2_1 _10282_ (.A(net589),
    .B(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__o32ai_1 _10283_ (.A1(_04928_),
    .A2(_04933_),
    .A3(_04937_),
    .B1(net540),
    .B2(\core.CPU_Xreg_value_a4[0][28] ),
    .Y(_04938_));
 sky130_fd_sc_hd__nor2_1 _10284_ (.A(_03457_),
    .B(net391),
    .Y(_04939_));
 sky130_fd_sc_hd__nor3_1 _10285_ (.A(_04625_),
    .B(_04939_),
    .C(net430),
    .Y(_04940_));
 sky130_fd_sc_hd__a21oi_1 _10286_ (.A1(net430),
    .A2(_04938_),
    .B1(_04940_),
    .Y(\core.CPU_src2_value_a2[28] ));
 sky130_fd_sc_hd__nand2b_1 _10287_ (.A_N(net587),
    .B(net592),
    .Y(_04941_));
 sky130_fd_sc_hd__mux2i_1 _10288_ (.A0(\core.CPU_Xreg_value_a4[1][29] ),
    .A1(\core.CPU_Xreg_value_a4[3][29] ),
    .S(net590),
    .Y(_04942_));
 sky130_fd_sc_hd__a21oi_1 _10289_ (.A1(_04164_),
    .A2(net590),
    .B1(net587),
    .Y(_04943_));
 sky130_fd_sc_hd__a21oi_1 _10290_ (.A1(\core.CPU_Xreg_value_a4[8][29] ),
    .A2(_04751_),
    .B1(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__mux2i_1 _10291_ (.A0(\core.CPU_Xreg_value_a4[10][29] ),
    .A1(\core.CPU_Xreg_value_a4[11][29] ),
    .S(\core.CPU_rf_rd_index2_a2[0] ),
    .Y(_04945_));
 sky130_fd_sc_hd__nand2_1 _10292_ (.A(\core.CPU_Xreg_value_a4[9][29] ),
    .B(net461),
    .Y(_04946_));
 sky130_fd_sc_hd__o21ai_0 _10293_ (.A1(net539),
    .A2(_04945_),
    .B1(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__nand2_1 _10294_ (.A(net587),
    .B(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__o221ai_1 _10295_ (.A1(_04941_),
    .A2(_04942_),
    .B1(_04944_),
    .B2(\core.CPU_rf_rd_index2_a2[0] ),
    .C1(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__o211ai_1 _10296_ (.A1(\core.CPU_Xreg_value_a4[0][29] ),
    .A2(net540),
    .B1(_04949_),
    .C1(net430),
    .Y(_04950_));
 sky130_fd_sc_hd__o31ai_1 _10297_ (.A1(_03506_),
    .A2(_03520_),
    .A3(net431),
    .B1(_04950_),
    .Y(\core.CPU_src2_value_a2[29] ));
 sky130_fd_sc_hd__mux4_2 _10298_ (.A0(\core.CPU_Xreg_value_a4[0][2] ),
    .A1(\core.CPU_Xreg_value_a4[1][2] ),
    .A2(\core.CPU_Xreg_value_a4[2][2] ),
    .A3(\core.CPU_Xreg_value_a4[3][2] ),
    .S0(net592),
    .S1(net590),
    .X(_04951_));
 sky130_fd_sc_hd__or3_1 _10299_ (.A(\core.CPU_Xreg_value_a4[0][2] ),
    .B(net587),
    .C(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__mux2_2 _10300_ (.A0(\core.CPU_Xreg_value_a4[10][2] ),
    .A1(\core.CPU_Xreg_value_a4[11][2] ),
    .S(net592),
    .X(_04953_));
 sky130_fd_sc_hd__nand2_1 _10301_ (.A(net590),
    .B(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__nand2_1 _10302_ (.A(\core.CPU_Xreg_value_a4[9][2] ),
    .B(net461),
    .Y(_04955_));
 sky130_fd_sc_hd__nor2_1 _10303_ (.A(net587),
    .B(_04951_),
    .Y(_04956_));
 sky130_fd_sc_hd__a31oi_1 _10304_ (.A1(net587),
    .A2(_04954_),
    .A3(_04955_),
    .B1(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__a31oi_2 _10305_ (.A1(\core.CPU_Xreg_value_a4[8][2] ),
    .A2(net537),
    .A3(_04952_),
    .B1(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__nor2_1 _10306_ (.A(\core.CPU_result_a3[2] ),
    .B(net431),
    .Y(_04959_));
 sky130_fd_sc_hd__a21oi_1 _10307_ (.A1(net431),
    .A2(_04958_),
    .B1(_04959_),
    .Y(\core.CPU_src2_value_a2[2] ));
 sky130_fd_sc_hd__mux4_2 _10308_ (.A0(\core.CPU_Xreg_value_a4[0][30] ),
    .A1(\core.CPU_Xreg_value_a4[1][30] ),
    .A2(\core.CPU_Xreg_value_a4[2][30] ),
    .A3(\core.CPU_Xreg_value_a4[3][30] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(\core.CPU_rf_rd_index2_a2[1] ),
    .X(_04960_));
 sky130_fd_sc_hd__mux4_2 _10309_ (.A0(\core.CPU_Xreg_value_a4[8][30] ),
    .A1(\core.CPU_Xreg_value_a4[9][30] ),
    .A2(\core.CPU_Xreg_value_a4[10][30] ),
    .A3(\core.CPU_Xreg_value_a4[11][30] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(\core.CPU_rf_rd_index2_a2[1] ),
    .X(_04961_));
 sky130_fd_sc_hd__mux2_2 _10310_ (.A0(_04960_),
    .A1(_04961_),
    .S(net588),
    .X(_04962_));
 sky130_fd_sc_hd__nand2_1 _10311_ (.A(net431),
    .B(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__o21ai_0 _10312_ (.A1(_04665_),
    .A2(net431),
    .B1(_04963_),
    .Y(\core.CPU_src2_value_a2[30] ));
 sky130_fd_sc_hd__mux2_2 _10313_ (.A0(\core.CPU_Xreg_value_a4[9][31] ),
    .A1(\core.CPU_Xreg_value_a4[11][31] ),
    .S(net590),
    .X(_04964_));
 sky130_fd_sc_hd__a22o_1 _10314_ (.A1(\core.CPU_Xreg_value_a4[3][31] ),
    .A2(net462),
    .B1(_04964_),
    .B2(net587),
    .X(_04965_));
 sky130_fd_sc_hd__o21ai_0 _10315_ (.A1(\core.CPU_Xreg_value_a4[2][31] ),
    .A2(_04751_),
    .B1(net538),
    .Y(_04966_));
 sky130_fd_sc_hd__a21boi_0 _10316_ (.A1(\core.CPU_Xreg_value_a4[1][31] ),
    .A2(_04751_),
    .B1_N(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__mux2i_1 _10317_ (.A0(\core.CPU_Xreg_value_a4[8][31] ),
    .A1(\core.CPU_Xreg_value_a4[10][31] ),
    .S(net590),
    .Y(_04968_));
 sky130_fd_sc_hd__o22ai_1 _10318_ (.A1(net587),
    .A2(_04967_),
    .B1(_04968_),
    .B2(_04831_),
    .Y(_04969_));
 sky130_fd_sc_hd__a21oi_1 _10319_ (.A1(\core.CPU_rf_rd_index2_a2[0] ),
    .A2(_04965_),
    .B1(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__nor2_1 _10320_ (.A(\core.CPU_Xreg_value_a4[0][31] ),
    .B(net540),
    .Y(_04971_));
 sky130_fd_sc_hd__o21ai_0 _10321_ (.A1(_04970_),
    .A2(_04971_),
    .B1(net430),
    .Y(_04972_));
 sky130_fd_sc_hd__o21a_1 _10322_ (.A1(_04673_),
    .A2(net430),
    .B1(_04972_),
    .X(\core.CPU_src2_value_a2[31] ));
 sky130_fd_sc_hd__a22o_1 _10323_ (.A1(\core.CPU_Xreg_value_a4[9][3] ),
    .A2(net461),
    .B1(net459),
    .B2(\core.CPU_Xreg_value_a4[10][3] ),
    .X(_04973_));
 sky130_fd_sc_hd__mux2i_1 _10324_ (.A0(\core.CPU_Xreg_value_a4[2][3] ),
    .A1(\core.CPU_Xreg_value_a4[3][3] ),
    .S(net592),
    .Y(_04974_));
 sky130_fd_sc_hd__nand3_1 _10325_ (.A(\core.CPU_Xreg_value_a4[11][3] ),
    .B(net587),
    .C(net592),
    .Y(_04975_));
 sky130_fd_sc_hd__o21ai_0 _10326_ (.A1(net587),
    .A2(_04974_),
    .B1(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__nor2_1 _10327_ (.A(\core.CPU_Xreg_value_a4[1][3] ),
    .B(net538),
    .Y(_04977_));
 sky130_fd_sc_hd__a2bb2oi_1 _10328_ (.A1_N(net587),
    .A2_N(_04977_),
    .B1(net538),
    .B2(\core.CPU_Xreg_value_a4[8][3] ),
    .Y(_04978_));
 sky130_fd_sc_hd__nor2_1 _10329_ (.A(net590),
    .B(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__a221o_1 _10330_ (.A1(net587),
    .A2(_04973_),
    .B1(_04976_),
    .B2(net590),
    .C1(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__o21ai_1 _10331_ (.A1(\core.CPU_Xreg_value_a4[0][3] ),
    .A2(net540),
    .B1(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__nor2_1 _10332_ (.A(net372),
    .B(net431),
    .Y(_04982_));
 sky130_fd_sc_hd__a21oi_1 _10333_ (.A1(net431),
    .A2(net385),
    .B1(_04982_),
    .Y(\core.CPU_src2_value_a2[3] ));
 sky130_fd_sc_hd__a22o_1 _10334_ (.A1(\core.CPU_Xreg_value_a4[9][4] ),
    .A2(_04760_),
    .B1(net459),
    .B2(\core.CPU_Xreg_value_a4[10][4] ),
    .X(_04983_));
 sky130_fd_sc_hd__mux2i_1 _10335_ (.A0(\core.CPU_Xreg_value_a4[2][4] ),
    .A1(\core.CPU_Xreg_value_a4[3][4] ),
    .S(net592),
    .Y(_04984_));
 sky130_fd_sc_hd__nand3_1 _10336_ (.A(\core.CPU_Xreg_value_a4[11][4] ),
    .B(net587),
    .C(net592),
    .Y(_04985_));
 sky130_fd_sc_hd__o21ai_0 _10337_ (.A1(net587),
    .A2(_04984_),
    .B1(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__inv_1 _10338_ (.A(\core.CPU_Xreg_value_a4[1][4] ),
    .Y(_04987_));
 sky130_fd_sc_hd__a21oi_1 _10339_ (.A1(_04987_),
    .A2(net592),
    .B1(net587),
    .Y(_04988_));
 sky130_fd_sc_hd__a21oi_1 _10340_ (.A1(\core.CPU_Xreg_value_a4[8][4] ),
    .A2(net538),
    .B1(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__nor2_1 _10341_ (.A(net590),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__a221o_1 _10342_ (.A1(net587),
    .A2(_04983_),
    .B1(_04986_),
    .B2(net590),
    .C1(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__o211ai_1 _10343_ (.A1(\core.CPU_Xreg_value_a4[0][4] ),
    .A2(net540),
    .B1(_04991_),
    .C1(net430),
    .Y(_04992_));
 sky130_fd_sc_hd__o21ai_0 _10344_ (.A1(_03659_),
    .A2(net431),
    .B1(net384),
    .Y(\core.CPU_src2_value_a2[4] ));
 sky130_fd_sc_hd__mux2i_1 _10345_ (.A0(\core.CPU_Xreg_value_a4[8][5] ),
    .A1(\core.CPU_Xreg_value_a4[9][5] ),
    .S(net592),
    .Y(_04993_));
 sky130_fd_sc_hd__nand2_1 _10346_ (.A(net587),
    .B(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__o21ai_0 _10347_ (.A1(\core.CPU_Xreg_value_a4[1][5] ),
    .A2(_04941_),
    .B1(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__mux4_2 _10348_ (.A0(\core.CPU_Xreg_value_a4[2][5] ),
    .A1(\core.CPU_Xreg_value_a4[3][5] ),
    .A2(\core.CPU_Xreg_value_a4[10][5] ),
    .A3(\core.CPU_Xreg_value_a4[11][5] ),
    .S0(net592),
    .S1(net587),
    .X(_04996_));
 sky130_fd_sc_hd__nand2_1 _10349_ (.A(net590),
    .B(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__o21ai_0 _10350_ (.A1(net590),
    .A2(_04995_),
    .B1(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__o211ai_1 _10351_ (.A1(\core.CPU_Xreg_value_a4[0][5] ),
    .A2(net540),
    .B1(_04998_),
    .C1(net430),
    .Y(_04999_));
 sky130_fd_sc_hd__o21ai_0 _10352_ (.A1(_03675_),
    .A2(net431),
    .B1(net395),
    .Y(\core.CPU_src2_value_a2[5] ));
 sky130_fd_sc_hd__mux4_2 _10353_ (.A0(\core.CPU_Xreg_value_a4[0][6] ),
    .A1(\core.CPU_Xreg_value_a4[1][6] ),
    .A2(\core.CPU_Xreg_value_a4[2][6] ),
    .A3(\core.CPU_Xreg_value_a4[3][6] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(\core.CPU_rf_rd_index2_a2[1] ),
    .X(_05000_));
 sky130_fd_sc_hd__mux4_2 _10354_ (.A0(\core.CPU_Xreg_value_a4[8][6] ),
    .A1(\core.CPU_Xreg_value_a4[9][6] ),
    .A2(\core.CPU_Xreg_value_a4[10][6] ),
    .A3(\core.CPU_Xreg_value_a4[11][6] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(\core.CPU_rf_rd_index2_a2[1] ),
    .X(_05001_));
 sky130_fd_sc_hd__mux2_2 _10355_ (.A0(_05000_),
    .A1(_05001_),
    .S(net587),
    .X(_05002_));
 sky130_fd_sc_hd__nand2_1 _10356_ (.A(net430),
    .B(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__o21ai_0 _10357_ (.A1(_03694_),
    .A2(net431),
    .B1(_05003_),
    .Y(\core.CPU_src2_value_a2[6] ));
 sky130_fd_sc_hd__mux4_2 _10358_ (.A0(\core.CPU_Xreg_value_a4[0][7] ),
    .A1(\core.CPU_Xreg_value_a4[1][7] ),
    .A2(\core.CPU_Xreg_value_a4[2][7] ),
    .A3(\core.CPU_Xreg_value_a4[3][7] ),
    .S0(net591),
    .S1(net589),
    .X(_05004_));
 sky130_fd_sc_hd__mux4_2 _10359_ (.A0(\core.CPU_Xreg_value_a4[8][7] ),
    .A1(\core.CPU_Xreg_value_a4[9][7] ),
    .A2(\core.CPU_Xreg_value_a4[10][7] ),
    .A3(\core.CPU_Xreg_value_a4[11][7] ),
    .S0(\core.CPU_rf_rd_index2_a2[0] ),
    .S1(\core.CPU_rf_rd_index2_a2[1] ),
    .X(_05005_));
 sky130_fd_sc_hd__mux2i_1 _10360_ (.A0(_05004_),
    .A1(_05005_),
    .S(net588),
    .Y(_05006_));
 sky130_fd_sc_hd__nor2_1 _10361_ (.A(_03706_),
    .B(net431),
    .Y(_05007_));
 sky130_fd_sc_hd__a21oi_1 _10362_ (.A1(net431),
    .A2(_05006_),
    .B1(_05007_),
    .Y(\core.CPU_src2_value_a2[7] ));
 sky130_fd_sc_hd__mux2_2 _10363_ (.A0(\core.CPU_Xreg_value_a4[9][8] ),
    .A1(\core.CPU_Xreg_value_a4[11][8] ),
    .S(net589),
    .X(_05008_));
 sky130_fd_sc_hd__a22oi_1 _10364_ (.A1(\core.CPU_Xreg_value_a4[3][8] ),
    .A2(net462),
    .B1(_05008_),
    .B2(\core.CPU_rf_rd_index2_a2[3] ),
    .Y(_05009_));
 sky130_fd_sc_hd__o21ai_0 _10365_ (.A1(\core.CPU_Xreg_value_a4[2][8] ),
    .A2(net539),
    .B1(net538),
    .Y(_05010_));
 sky130_fd_sc_hd__a21boi_0 _10366_ (.A1(\core.CPU_Xreg_value_a4[1][8] ),
    .A2(net539),
    .B1_N(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__mux2i_1 _10367_ (.A0(\core.CPU_Xreg_value_a4[8][8] ),
    .A1(\core.CPU_Xreg_value_a4[10][8] ),
    .S(net589),
    .Y(_05012_));
 sky130_fd_sc_hd__o22a_1 _10368_ (.A1(\core.CPU_rf_rd_index2_a2[3] ),
    .A2(_05011_),
    .B1(_05012_),
    .B2(_04831_),
    .X(_05013_));
 sky130_fd_sc_hd__o21ai_0 _10369_ (.A1(net538),
    .A2(_05009_),
    .B1(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__o21ai_0 _10370_ (.A1(\core.CPU_Xreg_value_a4[0][8] ),
    .A2(net540),
    .B1(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__nor2_1 _10371_ (.A(_04733_),
    .B(net431),
    .Y(_05016_));
 sky130_fd_sc_hd__a21oi_1 _10372_ (.A1(net431),
    .A2(net383),
    .B1(_05016_),
    .Y(\core.CPU_src2_value_a2[8] ));
 sky130_fd_sc_hd__a22o_1 _10373_ (.A1(\core.CPU_Xreg_value_a4[9][9] ),
    .A2(net461),
    .B1(_04816_),
    .B2(\core.CPU_Xreg_value_a4[10][9] ),
    .X(_05017_));
 sky130_fd_sc_hd__mux2i_1 _10374_ (.A0(\core.CPU_Xreg_value_a4[2][9] ),
    .A1(\core.CPU_Xreg_value_a4[3][9] ),
    .S(net591),
    .Y(_05018_));
 sky130_fd_sc_hd__nand3_1 _10375_ (.A(\core.CPU_Xreg_value_a4[11][9] ),
    .B(\core.CPU_rf_rd_index2_a2[3] ),
    .C(net591),
    .Y(_05019_));
 sky130_fd_sc_hd__o21ai_0 _10376_ (.A1(\core.CPU_rf_rd_index2_a2[3] ),
    .A2(_05018_),
    .B1(_05019_),
    .Y(_05020_));
 sky130_fd_sc_hd__nor2_1 _10377_ (.A(\core.CPU_Xreg_value_a4[1][9] ),
    .B(net538),
    .Y(_05021_));
 sky130_fd_sc_hd__a2bb2oi_1 _10378_ (.A1_N(\core.CPU_rf_rd_index2_a2[3] ),
    .A2_N(_05021_),
    .B1(net538),
    .B2(\core.CPU_Xreg_value_a4[8][9] ),
    .Y(_05022_));
 sky130_fd_sc_hd__nor2_1 _10379_ (.A(net589),
    .B(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__a221o_1 _10380_ (.A1(\core.CPU_rf_rd_index2_a2[3] ),
    .A2(_05017_),
    .B1(_05020_),
    .B2(net589),
    .C1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__o21ai_0 _10381_ (.A1(\core.CPU_Xreg_value_a4[0][9] ),
    .A2(_04748_),
    .B1(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__nor2_1 _10382_ (.A(_03741_),
    .B(net431),
    .Y(_05026_));
 sky130_fd_sc_hd__a21oi_1 _10383_ (.A1(net431),
    .A2(net382),
    .B1(_05026_),
    .Y(\core.CPU_src2_value_a2[9] ));
 sky130_fd_sc_hd__a21oi_1 _10387_ (.A1(\core.CPU_Dmem_value_a5[3][0] ),
    .A2(net505),
    .B1(net559),
    .Y(_05030_));
 sky130_fd_sc_hd__a22oi_1 _10390_ (.A1(\core.CPU_Dmem_value_a5[13][0] ),
    .A2(_01582_),
    .B1(_01660_),
    .B2(\core.CPU_Dmem_value_a5[14][0] ),
    .Y(_05033_));
 sky130_fd_sc_hd__a22oi_1 _10393_ (.A1(\core.CPU_Dmem_value_a5[15][0] ),
    .A2(_01734_),
    .B1(net507),
    .B2(\core.CPU_Dmem_value_a5[2][0] ),
    .Y(_05036_));
 sky130_fd_sc_hd__a22oi_1 _10396_ (.A1(\core.CPU_Dmem_value_a5[11][0] ),
    .A2(net528),
    .B1(net484),
    .B2(\core.CPU_Dmem_value_a5[8][0] ),
    .Y(_05039_));
 sky130_fd_sc_hd__nand4_1 _10397_ (.A(_05030_),
    .B(_05033_),
    .C(_05036_),
    .D(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__a22oi_1 _10400_ (.A1(\core.CPU_Dmem_value_a5[10][0] ),
    .A2(net530),
    .B1(net523),
    .B2(\core.CPU_Dmem_value_a5[12][0] ),
    .Y(_05043_));
 sky130_fd_sc_hd__a22oi_1 _10403_ (.A1(\core.CPU_Dmem_value_a5[1][0] ),
    .A2(net514),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][0] ),
    .Y(_05046_));
 sky130_fd_sc_hd__a22oi_1 _10406_ (.A1(\core.CPU_Dmem_value_a5[5][0] ),
    .A2(net498),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][0] ),
    .Y(_05049_));
 sky130_fd_sc_hd__a22oi_1 _10408_ (.A1(\core.CPU_Dmem_value_a5[7][0] ),
    .A2(_02275_),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][0] ),
    .Y(_05051_));
 sky130_fd_sc_hd__nand4_1 _10409_ (.A(_05043_),
    .B(_05046_),
    .C(_05049_),
    .D(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__o22a_1 _10410_ (.A1(\core.CPU_Dmem_value_a5[0][0] ),
    .A2(_01199_),
    .B1(_05040_),
    .B2(_05052_),
    .X(\core.w_CPU_dmem_rd_data_a4[0] ));
 sky130_fd_sc_hd__a21oi_1 _10411_ (.A1(\core.CPU_Dmem_value_a5[3][10] ),
    .A2(net505),
    .B1(net558),
    .Y(_05053_));
 sky130_fd_sc_hd__a22oi_1 _10414_ (.A1(\core.CPU_Dmem_value_a5[10][10] ),
    .A2(net530),
    .B1(net513),
    .B2(\core.CPU_Dmem_value_a5[1][10] ),
    .Y(_05056_));
 sky130_fd_sc_hd__a22oi_1 _10416_ (.A1(\core.CPU_Dmem_value_a5[14][10] ),
    .A2(net518),
    .B1(_02428_),
    .B2(\core.CPU_Dmem_value_a5[9][10] ),
    .Y(_05058_));
 sky130_fd_sc_hd__a22oi_1 _10418_ (.A1(\core.CPU_Dmem_value_a5[12][10] ),
    .A2(net524),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][10] ),
    .Y(_05060_));
 sky130_fd_sc_hd__nand4_1 _10419_ (.A(_05053_),
    .B(_05056_),
    .C(_05058_),
    .D(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__a22oi_1 _10422_ (.A1(\core.CPU_Dmem_value_a5[11][10] ),
    .A2(net527),
    .B1(net517),
    .B2(\core.CPU_Dmem_value_a5[15][10] ),
    .Y(_05064_));
 sky130_fd_sc_hd__a22oi_1 _10423_ (.A1(\core.CPU_Dmem_value_a5[2][10] ),
    .A2(net508),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][10] ),
    .Y(_05065_));
 sky130_fd_sc_hd__a22oi_1 _10426_ (.A1(\core.CPU_Dmem_value_a5[4][10] ),
    .A2(net499),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][10] ),
    .Y(_05068_));
 sky130_fd_sc_hd__a22oi_1 _10428_ (.A1(\core.CPU_Dmem_value_a5[5][10] ),
    .A2(net497),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][10] ),
    .Y(_05070_));
 sky130_fd_sc_hd__nand4_1 _10429_ (.A(_05064_),
    .B(_05065_),
    .C(_05068_),
    .D(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__o22a_1 _10430_ (.A1(\core.CPU_Dmem_value_a5[0][10] ),
    .A2(net534),
    .B1(_05061_),
    .B2(_05071_),
    .X(\core.w_CPU_dmem_rd_data_a4[10] ));
 sky130_fd_sc_hd__a21oi_1 _10432_ (.A1(\core.CPU_Dmem_value_a5[2][11] ),
    .A2(net508),
    .B1(net558),
    .Y(_05073_));
 sky130_fd_sc_hd__a22oi_1 _10434_ (.A1(\core.CPU_Dmem_value_a5[11][11] ),
    .A2(net527),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][11] ),
    .Y(_05075_));
 sky130_fd_sc_hd__a22oi_1 _10436_ (.A1(\core.CPU_Dmem_value_a5[14][11] ),
    .A2(net518),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][11] ),
    .Y(_05077_));
 sky130_fd_sc_hd__a22oi_1 _10437_ (.A1(\core.CPU_Dmem_value_a5[12][11] ),
    .A2(net524),
    .B1(net513),
    .B2(\core.CPU_Dmem_value_a5[1][11] ),
    .Y(_05078_));
 sky130_fd_sc_hd__nand4_1 _10438_ (.A(_05073_),
    .B(_05075_),
    .C(_05077_),
    .D(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__a22oi_1 _10439_ (.A1(\core.CPU_Dmem_value_a5[10][11] ),
    .A2(net529),
    .B1(net517),
    .B2(\core.CPU_Dmem_value_a5[15][11] ),
    .Y(_05080_));
 sky130_fd_sc_hd__a22oi_1 _10442_ (.A1(\core.CPU_Dmem_value_a5[3][11] ),
    .A2(net505),
    .B1(_02428_),
    .B2(\core.CPU_Dmem_value_a5[9][11] ),
    .Y(_05083_));
 sky130_fd_sc_hd__a22oi_1 _10444_ (.A1(\core.CPU_Dmem_value_a5[13][11] ),
    .A2(net522),
    .B1(net491),
    .B2(\core.CPU_Dmem_value_a5[6][11] ),
    .Y(_05085_));
 sky130_fd_sc_hd__a22oi_1 _10446_ (.A1(\core.CPU_Dmem_value_a5[4][11] ),
    .A2(net499),
    .B1(net497),
    .B2(\core.CPU_Dmem_value_a5[5][11] ),
    .Y(_05087_));
 sky130_fd_sc_hd__nand4_1 _10447_ (.A(_05080_),
    .B(_05083_),
    .C(_05085_),
    .D(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__o22a_1 _10448_ (.A1(\core.CPU_Dmem_value_a5[0][11] ),
    .A2(net534),
    .B1(_05079_),
    .B2(_05088_),
    .X(\core.w_CPU_dmem_rd_data_a4[11] ));
 sky130_fd_sc_hd__a21oi_1 _10450_ (.A1(\core.CPU_Dmem_value_a5[8][12] ),
    .A2(net485),
    .B1(net558),
    .Y(_05090_));
 sky130_fd_sc_hd__a22oi_1 _10452_ (.A1(\core.CPU_Dmem_value_a5[10][12] ),
    .A2(net529),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][12] ),
    .Y(_05092_));
 sky130_fd_sc_hd__a22oi_1 _10453_ (.A1(\core.CPU_Dmem_value_a5[14][12] ),
    .A2(net518),
    .B1(net491),
    .B2(\core.CPU_Dmem_value_a5[6][12] ),
    .Y(_05093_));
 sky130_fd_sc_hd__a22oi_1 _10455_ (.A1(\core.CPU_Dmem_value_a5[11][12] ),
    .A2(net527),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][12] ),
    .Y(_05095_));
 sky130_fd_sc_hd__nand4_1 _10456_ (.A(_05090_),
    .B(_05092_),
    .C(_05093_),
    .D(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__a22o_1 _10458_ (.A1(\core.CPU_Dmem_value_a5[2][12] ),
    .A2(net508),
    .B1(net505),
    .B2(\core.CPU_Dmem_value_a5[3][12] ),
    .X(_05098_));
 sky130_fd_sc_hd__a221oi_1 _10459_ (.A1(\core.CPU_Dmem_value_a5[1][12] ),
    .A2(net513),
    .B1(net497),
    .B2(\core.CPU_Dmem_value_a5[5][12] ),
    .C1(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__a22oi_1 _10460_ (.A1(\core.CPU_Dmem_value_a5[12][12] ),
    .A2(net524),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][12] ),
    .Y(_05100_));
 sky130_fd_sc_hd__a22oi_1 _10462_ (.A1(\core.CPU_Dmem_value_a5[15][12] ),
    .A2(net517),
    .B1(net499),
    .B2(\core.CPU_Dmem_value_a5[4][12] ),
    .Y(_05102_));
 sky130_fd_sc_hd__nand3_1 _10463_ (.A(_05099_),
    .B(_05100_),
    .C(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__o22a_1 _10464_ (.A1(\core.CPU_Dmem_value_a5[0][12] ),
    .A2(net534),
    .B1(_05096_),
    .B2(_05103_),
    .X(\core.w_CPU_dmem_rd_data_a4[12] ));
 sky130_fd_sc_hd__a21oi_1 _10465_ (.A1(\core.CPU_Dmem_value_a5[1][13] ),
    .A2(net514),
    .B1(net559),
    .Y(_05104_));
 sky130_fd_sc_hd__a22oi_1 _10466_ (.A1(\core.CPU_Dmem_value_a5[10][13] ),
    .A2(net530),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][13] ),
    .Y(_05105_));
 sky130_fd_sc_hd__a22oi_1 _10467_ (.A1(\core.CPU_Dmem_value_a5[14][13] ),
    .A2(_01660_),
    .B1(net506),
    .B2(\core.CPU_Dmem_value_a5[3][13] ),
    .Y(_05106_));
 sky130_fd_sc_hd__a22oi_1 _10468_ (.A1(\core.CPU_Dmem_value_a5[11][13] ),
    .A2(net528),
    .B1(_01734_),
    .B2(\core.CPU_Dmem_value_a5[15][13] ),
    .Y(_05107_));
 sky130_fd_sc_hd__nand4_1 _10469_ (.A(_05104_),
    .B(_05105_),
    .C(_05106_),
    .D(_05107_),
    .Y(_05108_));
 sky130_fd_sc_hd__a22oi_1 _10470_ (.A1(\core.CPU_Dmem_value_a5[12][13] ),
    .A2(net523),
    .B1(_01582_),
    .B2(\core.CPU_Dmem_value_a5[13][13] ),
    .Y(_05109_));
 sky130_fd_sc_hd__a22oi_1 _10471_ (.A1(\core.CPU_Dmem_value_a5[2][13] ),
    .A2(net507),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][13] ),
    .Y(_05110_));
 sky130_fd_sc_hd__a22oi_1 _10472_ (.A1(\core.CPU_Dmem_value_a5[8][13] ),
    .A2(net484),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][13] ),
    .Y(_05111_));
 sky130_fd_sc_hd__a22oi_1 _10474_ (.A1(\core.CPU_Dmem_value_a5[6][13] ),
    .A2(net492),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][13] ),
    .Y(_05113_));
 sky130_fd_sc_hd__nand4_1 _10475_ (.A(_05109_),
    .B(_05110_),
    .C(_05111_),
    .D(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__o22a_1 _10476_ (.A1(\core.CPU_Dmem_value_a5[0][13] ),
    .A2(_01199_),
    .B1(_05108_),
    .B2(_05114_),
    .X(\core.w_CPU_dmem_rd_data_a4[13] ));
 sky130_fd_sc_hd__a21oi_1 _10477_ (.A1(\core.CPU_Dmem_value_a5[9][14] ),
    .A2(net483),
    .B1(net558),
    .Y(_05115_));
 sky130_fd_sc_hd__a22oi_1 _10478_ (.A1(\core.CPU_Dmem_value_a5[10][14] ),
    .A2(net529),
    .B1(net524),
    .B2(\core.CPU_Dmem_value_a5[12][14] ),
    .Y(_05116_));
 sky130_fd_sc_hd__a22oi_1 _10479_ (.A1(\core.CPU_Dmem_value_a5[15][14] ),
    .A2(net517),
    .B1(net505),
    .B2(\core.CPU_Dmem_value_a5[3][14] ),
    .Y(_05117_));
 sky130_fd_sc_hd__a22oi_1 _10480_ (.A1(\core.CPU_Dmem_value_a5[11][14] ),
    .A2(net527),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][14] ),
    .Y(_05118_));
 sky130_fd_sc_hd__nand4_1 _10481_ (.A(_05115_),
    .B(_05116_),
    .C(_05117_),
    .D(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__a22o_1 _10482_ (.A1(\core.CPU_Dmem_value_a5[2][14] ),
    .A2(net508),
    .B1(_02275_),
    .B2(\core.CPU_Dmem_value_a5[7][14] ),
    .X(_05120_));
 sky130_fd_sc_hd__a221oi_1 _10483_ (.A1(\core.CPU_Dmem_value_a5[14][14] ),
    .A2(net518),
    .B1(net513),
    .B2(\core.CPU_Dmem_value_a5[1][14] ),
    .C1(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__a22oi_1 _10484_ (.A1(\core.CPU_Dmem_value_a5[5][14] ),
    .A2(net497),
    .B1(net491),
    .B2(\core.CPU_Dmem_value_a5[6][14] ),
    .Y(_05122_));
 sky130_fd_sc_hd__a22oi_1 _10485_ (.A1(\core.CPU_Dmem_value_a5[4][14] ),
    .A2(net499),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][14] ),
    .Y(_05123_));
 sky130_fd_sc_hd__nand3_1 _10486_ (.A(_05121_),
    .B(_05122_),
    .C(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__o22a_1 _10487_ (.A1(\core.CPU_Dmem_value_a5[0][14] ),
    .A2(net534),
    .B1(_05119_),
    .B2(_05124_),
    .X(\core.w_CPU_dmem_rd_data_a4[14] ));
 sky130_fd_sc_hd__a21oi_1 _10488_ (.A1(\core.CPU_Dmem_value_a5[8][15] ),
    .A2(net485),
    .B1(net559),
    .Y(_05125_));
 sky130_fd_sc_hd__a22oi_1 _10489_ (.A1(\core.CPU_Dmem_value_a5[11][15] ),
    .A2(net528),
    .B1(net518),
    .B2(\core.CPU_Dmem_value_a5[14][15] ),
    .Y(_05126_));
 sky130_fd_sc_hd__a22oi_1 _10490_ (.A1(\core.CPU_Dmem_value_a5[2][15] ),
    .A2(net508),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][15] ),
    .Y(_05127_));
 sky130_fd_sc_hd__a22oi_1 _10491_ (.A1(\core.CPU_Dmem_value_a5[12][15] ),
    .A2(net524),
    .B1(_02428_),
    .B2(\core.CPU_Dmem_value_a5[9][15] ),
    .Y(_05128_));
 sky130_fd_sc_hd__nand4_1 _10492_ (.A(_05125_),
    .B(_05126_),
    .C(_05127_),
    .D(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__a22oi_1 _10493_ (.A1(\core.CPU_Dmem_value_a5[10][15] ),
    .A2(net530),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][15] ),
    .Y(_05130_));
 sky130_fd_sc_hd__a22oi_1 _10494_ (.A1(\core.CPU_Dmem_value_a5[3][15] ),
    .A2(net506),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][15] ),
    .Y(_05131_));
 sky130_fd_sc_hd__a22oi_1 _10495_ (.A1(\core.CPU_Dmem_value_a5[13][15] ),
    .A2(net522),
    .B1(net514),
    .B2(\core.CPU_Dmem_value_a5[1][15] ),
    .Y(_05132_));
 sky130_fd_sc_hd__a22oi_1 _10496_ (.A1(\core.CPU_Dmem_value_a5[15][15] ),
    .A2(net517),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][15] ),
    .Y(_05133_));
 sky130_fd_sc_hd__nand4_1 _10497_ (.A(_05130_),
    .B(_05131_),
    .C(_05132_),
    .D(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__o22a_1 _10498_ (.A1(\core.CPU_Dmem_value_a5[0][15] ),
    .A2(net534),
    .B1(_05129_),
    .B2(_05134_),
    .X(\core.w_CPU_dmem_rd_data_a4[15] ));
 sky130_fd_sc_hd__a21oi_1 _10499_ (.A1(\core.CPU_Dmem_value_a5[3][16] ),
    .A2(net506),
    .B1(net559),
    .Y(_05135_));
 sky130_fd_sc_hd__a22oi_1 _10501_ (.A1(\core.CPU_Dmem_value_a5[12][16] ),
    .A2(net523),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][16] ),
    .Y(_05137_));
 sky130_fd_sc_hd__a22oi_1 _10502_ (.A1(\core.CPU_Dmem_value_a5[15][16] ),
    .A2(_01734_),
    .B1(net514),
    .B2(\core.CPU_Dmem_value_a5[1][16] ),
    .Y(_05138_));
 sky130_fd_sc_hd__a22oi_1 _10504_ (.A1(\core.CPU_Dmem_value_a5[13][16] ),
    .A2(_01582_),
    .B1(_01660_),
    .B2(\core.CPU_Dmem_value_a5[14][16] ),
    .Y(_05140_));
 sky130_fd_sc_hd__nand4_1 _10505_ (.A(_05135_),
    .B(_05137_),
    .C(_05138_),
    .D(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__a22oi_1 _10506_ (.A1(\core.CPU_Dmem_value_a5[10][16] ),
    .A2(net530),
    .B1(net528),
    .B2(\core.CPU_Dmem_value_a5[11][16] ),
    .Y(_05142_));
 sky130_fd_sc_hd__a22oi_1 _10507_ (.A1(\core.CPU_Dmem_value_a5[2][16] ),
    .A2(net507),
    .B1(net484),
    .B2(\core.CPU_Dmem_value_a5[8][16] ),
    .Y(_05143_));
 sky130_fd_sc_hd__a22oi_1 _10508_ (.A1(\core.CPU_Dmem_value_a5[5][16] ),
    .A2(net498),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][16] ),
    .Y(_05144_));
 sky130_fd_sc_hd__a22oi_1 _10509_ (.A1(\core.CPU_Dmem_value_a5[4][16] ),
    .A2(net500),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][16] ),
    .Y(_05145_));
 sky130_fd_sc_hd__nand4_1 _10510_ (.A(_05142_),
    .B(_05143_),
    .C(_05144_),
    .D(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__o22a_1 _10511_ (.A1(\core.CPU_Dmem_value_a5[0][16] ),
    .A2(_01199_),
    .B1(_05141_),
    .B2(_05146_),
    .X(\core.w_CPU_dmem_rd_data_a4[16] ));
 sky130_fd_sc_hd__a21oi_1 _10513_ (.A1(\core.CPU_Dmem_value_a5[7][17] ),
    .A2(net490),
    .B1(net559),
    .Y(_05148_));
 sky130_fd_sc_hd__a22oi_1 _10514_ (.A1(\core.CPU_Dmem_value_a5[13][17] ),
    .A2(_01582_),
    .B1(_01734_),
    .B2(\core.CPU_Dmem_value_a5[15][17] ),
    .Y(_05149_));
 sky130_fd_sc_hd__a22oi_1 _10515_ (.A1(\core.CPU_Dmem_value_a5[4][17] ),
    .A2(net500),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][17] ),
    .Y(_05150_));
 sky130_fd_sc_hd__a22oi_1 _10516_ (.A1(\core.CPU_Dmem_value_a5[12][17] ),
    .A2(net523),
    .B1(_01660_),
    .B2(\core.CPU_Dmem_value_a5[14][17] ),
    .Y(_05151_));
 sky130_fd_sc_hd__nand4_1 _10517_ (.A(_05148_),
    .B(_05149_),
    .C(_05150_),
    .D(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__a22o_1 _10518_ (.A1(\core.CPU_Dmem_value_a5[3][17] ),
    .A2(net506),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][17] ),
    .X(_05153_));
 sky130_fd_sc_hd__a221oi_1 _10519_ (.A1(\core.CPU_Dmem_value_a5[1][17] ),
    .A2(net514),
    .B1(net507),
    .B2(\core.CPU_Dmem_value_a5[2][17] ),
    .C1(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__a22oi_1 _10520_ (.A1(\core.CPU_Dmem_value_a5[11][17] ),
    .A2(net528),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][17] ),
    .Y(_05155_));
 sky130_fd_sc_hd__a22oi_1 _10521_ (.A1(\core.CPU_Dmem_value_a5[10][17] ),
    .A2(net530),
    .B1(net484),
    .B2(\core.CPU_Dmem_value_a5[8][17] ),
    .Y(_05156_));
 sky130_fd_sc_hd__nand3_1 _10522_ (.A(_05154_),
    .B(_05155_),
    .C(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__o22a_1 _10523_ (.A1(\core.CPU_Dmem_value_a5[0][17] ),
    .A2(_01199_),
    .B1(_05152_),
    .B2(_05157_),
    .X(\core.w_CPU_dmem_rd_data_a4[17] ));
 sky130_fd_sc_hd__a21oi_1 _10524_ (.A1(\core.CPU_Dmem_value_a5[8][18] ),
    .A2(net484),
    .B1(net559),
    .Y(_05158_));
 sky130_fd_sc_hd__a22oi_1 _10525_ (.A1(\core.CPU_Dmem_value_a5[13][18] ),
    .A2(_01582_),
    .B1(_01734_),
    .B2(\core.CPU_Dmem_value_a5[15][18] ),
    .Y(_05159_));
 sky130_fd_sc_hd__a22oi_1 _10526_ (.A1(\core.CPU_Dmem_value_a5[4][18] ),
    .A2(net500),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][18] ),
    .Y(_05160_));
 sky130_fd_sc_hd__a22oi_1 _10527_ (.A1(\core.CPU_Dmem_value_a5[11][18] ),
    .A2(net528),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][18] ),
    .Y(_05161_));
 sky130_fd_sc_hd__nand4_1 _10528_ (.A(_05158_),
    .B(_05159_),
    .C(_05160_),
    .D(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__a22oi_1 _10529_ (.A1(\core.CPU_Dmem_value_a5[10][18] ),
    .A2(net530),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][18] ),
    .Y(_05163_));
 sky130_fd_sc_hd__a22oi_1 _10530_ (.A1(\core.CPU_Dmem_value_a5[1][18] ),
    .A2(net514),
    .B1(net507),
    .B2(\core.CPU_Dmem_value_a5[2][18] ),
    .Y(_05164_));
 sky130_fd_sc_hd__a22oi_1 _10531_ (.A1(\core.CPU_Dmem_value_a5[12][18] ),
    .A2(net523),
    .B1(net506),
    .B2(\core.CPU_Dmem_value_a5[3][18] ),
    .Y(_05165_));
 sky130_fd_sc_hd__a22oi_1 _10532_ (.A1(\core.CPU_Dmem_value_a5[14][18] ),
    .A2(_01660_),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][18] ),
    .Y(_05166_));
 sky130_fd_sc_hd__nand4_1 _10533_ (.A(_05163_),
    .B(_05164_),
    .C(_05165_),
    .D(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__o22a_1 _10534_ (.A1(\core.CPU_Dmem_value_a5[0][18] ),
    .A2(_01199_),
    .B1(_05162_),
    .B2(_05167_),
    .X(\core.w_CPU_dmem_rd_data_a4[18] ));
 sky130_fd_sc_hd__a21oi_1 _10536_ (.A1(\core.CPU_Dmem_value_a5[8][19] ),
    .A2(net485),
    .B1(net558),
    .Y(_05169_));
 sky130_fd_sc_hd__a22oi_1 _10537_ (.A1(\core.CPU_Dmem_value_a5[12][19] ),
    .A2(net524),
    .B1(net513),
    .B2(\core.CPU_Dmem_value_a5[1][19] ),
    .Y(_05170_));
 sky130_fd_sc_hd__a22oi_1 _10538_ (.A1(\core.CPU_Dmem_value_a5[13][19] ),
    .A2(net522),
    .B1(net491),
    .B2(\core.CPU_Dmem_value_a5[6][19] ),
    .Y(_05171_));
 sky130_fd_sc_hd__a22oi_1 _10540_ (.A1(\core.CPU_Dmem_value_a5[10][19] ),
    .A2(net529),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][19] ),
    .Y(_05173_));
 sky130_fd_sc_hd__nand4_1 _10541_ (.A(_05169_),
    .B(_05170_),
    .C(_05171_),
    .D(_05173_),
    .Y(_05174_));
 sky130_fd_sc_hd__a22o_1 _10542_ (.A1(\core.CPU_Dmem_value_a5[2][19] ),
    .A2(net508),
    .B1(_02428_),
    .B2(\core.CPU_Dmem_value_a5[9][19] ),
    .X(_05175_));
 sky130_fd_sc_hd__a221oi_1 _10543_ (.A1(\core.CPU_Dmem_value_a5[14][19] ),
    .A2(net518),
    .B1(net505),
    .B2(\core.CPU_Dmem_value_a5[3][19] ),
    .C1(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__a22oi_1 _10544_ (.A1(\core.CPU_Dmem_value_a5[11][19] ),
    .A2(net527),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][19] ),
    .Y(_05177_));
 sky130_fd_sc_hd__a22oi_1 _10545_ (.A1(\core.CPU_Dmem_value_a5[15][19] ),
    .A2(net517),
    .B1(net497),
    .B2(\core.CPU_Dmem_value_a5[5][19] ),
    .Y(_05178_));
 sky130_fd_sc_hd__nand3_1 _10546_ (.A(_05176_),
    .B(_05177_),
    .C(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__o22a_1 _10547_ (.A1(\core.CPU_Dmem_value_a5[0][19] ),
    .A2(net534),
    .B1(_05174_),
    .B2(_05179_),
    .X(\core.w_CPU_dmem_rd_data_a4[19] ));
 sky130_fd_sc_hd__a22oi_1 _10548_ (.A1(\core.CPU_Dmem_value_a5[12][1] ),
    .A2(net523),
    .B1(_01660_),
    .B2(\core.CPU_Dmem_value_a5[14][1] ),
    .Y(_05180_));
 sky130_fd_sc_hd__a22oi_1 _10549_ (.A1(\core.CPU_Dmem_value_a5[11][1] ),
    .A2(net528),
    .B1(net506),
    .B2(\core.CPU_Dmem_value_a5[3][1] ),
    .Y(_05181_));
 sky130_fd_sc_hd__a22oi_1 _10551_ (.A1(\core.CPU_Dmem_value_a5[15][1] ),
    .A2(_01734_),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][1] ),
    .Y(_05183_));
 sky130_fd_sc_hd__a22oi_1 _10552_ (.A1(\core.CPU_Dmem_value_a5[10][1] ),
    .A2(net530),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][1] ),
    .Y(_05184_));
 sky130_fd_sc_hd__nand4_1 _10553_ (.A(_05180_),
    .B(_05181_),
    .C(_05183_),
    .D(_05184_),
    .Y(_05185_));
 sky130_fd_sc_hd__a22oi_1 _10554_ (.A1(\core.CPU_Dmem_value_a5[13][1] ),
    .A2(net522),
    .B1(net508),
    .B2(\core.CPU_Dmem_value_a5[2][1] ),
    .Y(_05186_));
 sky130_fd_sc_hd__a22oi_1 _10555_ (.A1(\core.CPU_Dmem_value_a5[1][1] ),
    .A2(net514),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][1] ),
    .Y(_05187_));
 sky130_fd_sc_hd__a22oi_1 _10556_ (.A1(\core.CPU_Dmem_value_a5[6][1] ),
    .A2(net492),
    .B1(net484),
    .B2(\core.CPU_Dmem_value_a5[8][1] ),
    .Y(_05188_));
 sky130_fd_sc_hd__a21oi_1 _10558_ (.A1(\core.CPU_Dmem_value_a5[9][1] ),
    .A2(net483),
    .B1(net559),
    .Y(_05190_));
 sky130_fd_sc_hd__nand4_1 _10559_ (.A(_05186_),
    .B(_05187_),
    .C(_05188_),
    .D(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__o22a_1 _10560_ (.A1(\core.CPU_Dmem_value_a5[0][1] ),
    .A2(net534),
    .B1(_05185_),
    .B2(_05191_),
    .X(\core.w_CPU_dmem_rd_data_a4[1] ));
 sky130_fd_sc_hd__a21oi_1 _10561_ (.A1(\core.CPU_Dmem_value_a5[2][20] ),
    .A2(net508),
    .B1(net559),
    .Y(_05192_));
 sky130_fd_sc_hd__a22oi_1 _10562_ (.A1(\core.CPU_Dmem_value_a5[10][20] ),
    .A2(net530),
    .B1(net497),
    .B2(\core.CPU_Dmem_value_a5[5][20] ),
    .Y(_05193_));
 sky130_fd_sc_hd__a22oi_1 _10563_ (.A1(\core.CPU_Dmem_value_a5[4][20] ),
    .A2(net500),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][20] ),
    .Y(_05194_));
 sky130_fd_sc_hd__a22oi_1 _10564_ (.A1(\core.CPU_Dmem_value_a5[11][20] ),
    .A2(net528),
    .B1(net518),
    .B2(\core.CPU_Dmem_value_a5[14][20] ),
    .Y(_05195_));
 sky130_fd_sc_hd__nand4_1 _10565_ (.A(_05192_),
    .B(_05193_),
    .C(_05194_),
    .D(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__a22oi_1 _10566_ (.A1(\core.CPU_Dmem_value_a5[12][20] ),
    .A2(net524),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][20] ),
    .Y(_05197_));
 sky130_fd_sc_hd__a22oi_1 _10567_ (.A1(\core.CPU_Dmem_value_a5[1][20] ),
    .A2(net514),
    .B1(net505),
    .B2(\core.CPU_Dmem_value_a5[3][20] ),
    .Y(_05198_));
 sky130_fd_sc_hd__a22oi_1 _10568_ (.A1(\core.CPU_Dmem_value_a5[15][20] ),
    .A2(net517),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][20] ),
    .Y(_05199_));
 sky130_fd_sc_hd__a22oi_1 _10569_ (.A1(\core.CPU_Dmem_value_a5[7][20] ),
    .A2(net490),
    .B1(_02428_),
    .B2(\core.CPU_Dmem_value_a5[9][20] ),
    .Y(_05200_));
 sky130_fd_sc_hd__nand4_1 _10570_ (.A(_05197_),
    .B(_05198_),
    .C(_05199_),
    .D(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__o22a_1 _10571_ (.A1(\core.CPU_Dmem_value_a5[0][20] ),
    .A2(net534),
    .B1(_05196_),
    .B2(_05201_),
    .X(\core.w_CPU_dmem_rd_data_a4[20] ));
 sky130_fd_sc_hd__a21oi_1 _10572_ (.A1(\core.CPU_Dmem_value_a5[9][21] ),
    .A2(_02428_),
    .B1(net559),
    .Y(_05202_));
 sky130_fd_sc_hd__a22oi_1 _10573_ (.A1(\core.CPU_Dmem_value_a5[10][21] ),
    .A2(net530),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][21] ),
    .Y(_05203_));
 sky130_fd_sc_hd__a22oi_1 _10574_ (.A1(\core.CPU_Dmem_value_a5[5][21] ),
    .A2(net498),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][21] ),
    .Y(_05204_));
 sky130_fd_sc_hd__a22oi_1 _10575_ (.A1(\core.CPU_Dmem_value_a5[14][21] ),
    .A2(net518),
    .B1(net517),
    .B2(\core.CPU_Dmem_value_a5[15][21] ),
    .Y(_05205_));
 sky130_fd_sc_hd__nand4_1 _10576_ (.A(_05202_),
    .B(_05203_),
    .C(_05204_),
    .D(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__a22o_1 _10577_ (.A1(\core.CPU_Dmem_value_a5[3][21] ),
    .A2(net506),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][21] ),
    .X(_05207_));
 sky130_fd_sc_hd__a221oi_1 _10578_ (.A1(\core.CPU_Dmem_value_a5[12][21] ),
    .A2(net524),
    .B1(net507),
    .B2(\core.CPU_Dmem_value_a5[2][21] ),
    .C1(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__a22oi_1 _10579_ (.A1(\core.CPU_Dmem_value_a5[11][21] ),
    .A2(net528),
    .B1(net514),
    .B2(\core.CPU_Dmem_value_a5[1][21] ),
    .Y(_05209_));
 sky130_fd_sc_hd__a22oi_1 _10580_ (.A1(\core.CPU_Dmem_value_a5[13][21] ),
    .A2(net522),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][21] ),
    .Y(_05210_));
 sky130_fd_sc_hd__nand3_1 _10581_ (.A(_05208_),
    .B(_05209_),
    .C(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__o22a_1 _10582_ (.A1(\core.CPU_Dmem_value_a5[0][21] ),
    .A2(net534),
    .B1(_05206_),
    .B2(_05211_),
    .X(\core.w_CPU_dmem_rd_data_a4[21] ));
 sky130_fd_sc_hd__a22oi_1 _10583_ (.A1(\core.CPU_Dmem_value_a5[12][22] ),
    .A2(net524),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][22] ),
    .Y(_05212_));
 sky130_fd_sc_hd__a22oi_1 _10584_ (.A1(\core.CPU_Dmem_value_a5[10][22] ),
    .A2(net530),
    .B1(net499),
    .B2(\core.CPU_Dmem_value_a5[4][22] ),
    .Y(_05213_));
 sky130_fd_sc_hd__a22oi_1 _10585_ (.A1(\core.CPU_Dmem_value_a5[14][22] ),
    .A2(net518),
    .B1(net513),
    .B2(\core.CPU_Dmem_value_a5[1][22] ),
    .Y(_05214_));
 sky130_fd_sc_hd__a22oi_1 _10586_ (.A1(\core.CPU_Dmem_value_a5[11][22] ),
    .A2(net527),
    .B1(_02428_),
    .B2(\core.CPU_Dmem_value_a5[9][22] ),
    .Y(_05215_));
 sky130_fd_sc_hd__nand4_1 _10587_ (.A(_05212_),
    .B(_05213_),
    .C(_05214_),
    .D(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__a22oi_1 _10588_ (.A1(\core.CPU_Dmem_value_a5[15][22] ),
    .A2(net517),
    .B1(net508),
    .B2(\core.CPU_Dmem_value_a5[2][22] ),
    .Y(_05217_));
 sky130_fd_sc_hd__a22oi_1 _10589_ (.A1(\core.CPU_Dmem_value_a5[3][22] ),
    .A2(net505),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][22] ),
    .Y(_05218_));
 sky130_fd_sc_hd__a22oi_1 _10590_ (.A1(\core.CPU_Dmem_value_a5[5][22] ),
    .A2(net497),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][22] ),
    .Y(_05219_));
 sky130_fd_sc_hd__a21oi_1 _10591_ (.A1(\core.CPU_Dmem_value_a5[8][22] ),
    .A2(net485),
    .B1(net558),
    .Y(_05220_));
 sky130_fd_sc_hd__nand4_1 _10592_ (.A(_05217_),
    .B(_05218_),
    .C(_05219_),
    .D(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__o22a_1 _10593_ (.A1(\core.CPU_Dmem_value_a5[0][22] ),
    .A2(net534),
    .B1(_05216_),
    .B2(_05221_),
    .X(\core.w_CPU_dmem_rd_data_a4[22] ));
 sky130_fd_sc_hd__a21oi_1 _10594_ (.A1(\core.CPU_Dmem_value_a5[2][23] ),
    .A2(net508),
    .B1(net558),
    .Y(_05222_));
 sky130_fd_sc_hd__a22oi_1 _10595_ (.A1(\core.CPU_Dmem_value_a5[10][23] ),
    .A2(net530),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][23] ),
    .Y(_05223_));
 sky130_fd_sc_hd__a22oi_1 _10596_ (.A1(\core.CPU_Dmem_value_a5[11][23] ),
    .A2(net527),
    .B1(net513),
    .B2(\core.CPU_Dmem_value_a5[1][23] ),
    .Y(_05224_));
 sky130_fd_sc_hd__a22oi_1 _10597_ (.A1(\core.CPU_Dmem_value_a5[13][23] ),
    .A2(net522),
    .B1(net518),
    .B2(\core.CPU_Dmem_value_a5[14][23] ),
    .Y(_05225_));
 sky130_fd_sc_hd__nand4_1 _10598_ (.A(_05222_),
    .B(_05223_),
    .C(_05224_),
    .D(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__a22oi_1 _10599_ (.A1(\core.CPU_Dmem_value_a5[12][23] ),
    .A2(net524),
    .B1(net517),
    .B2(\core.CPU_Dmem_value_a5[15][23] ),
    .Y(_05227_));
 sky130_fd_sc_hd__a22oi_1 _10600_ (.A1(\core.CPU_Dmem_value_a5[3][23] ),
    .A2(net505),
    .B1(net497),
    .B2(\core.CPU_Dmem_value_a5[5][23] ),
    .Y(_05228_));
 sky130_fd_sc_hd__a22oi_1 _10601_ (.A1(\core.CPU_Dmem_value_a5[4][23] ),
    .A2(net499),
    .B1(net491),
    .B2(\core.CPU_Dmem_value_a5[6][23] ),
    .Y(_05229_));
 sky130_fd_sc_hd__a22oi_1 _10602_ (.A1(\core.CPU_Dmem_value_a5[7][23] ),
    .A2(net490),
    .B1(_02428_),
    .B2(\core.CPU_Dmem_value_a5[9][23] ),
    .Y(_05230_));
 sky130_fd_sc_hd__nand4_1 _10603_ (.A(_05227_),
    .B(_05228_),
    .C(_05229_),
    .D(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__o22a_1 _10604_ (.A1(\core.CPU_Dmem_value_a5[0][23] ),
    .A2(net534),
    .B1(_05226_),
    .B2(_05231_),
    .X(\core.w_CPU_dmem_rd_data_a4[23] ));
 sky130_fd_sc_hd__a22oi_1 _10605_ (.A1(\core.CPU_Dmem_value_a5[10][24] ),
    .A2(net530),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][24] ),
    .Y(_05232_));
 sky130_fd_sc_hd__a22oi_1 _10606_ (.A1(\core.CPU_Dmem_value_a5[14][24] ),
    .A2(net518),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][24] ),
    .Y(_05233_));
 sky130_fd_sc_hd__a22oi_1 _10607_ (.A1(\core.CPU_Dmem_value_a5[15][24] ),
    .A2(net517),
    .B1(net514),
    .B2(\core.CPU_Dmem_value_a5[1][24] ),
    .Y(_05234_));
 sky130_fd_sc_hd__a22oi_1 _10608_ (.A1(\core.CPU_Dmem_value_a5[11][24] ),
    .A2(net527),
    .B1(net497),
    .B2(\core.CPU_Dmem_value_a5[5][24] ),
    .Y(_05235_));
 sky130_fd_sc_hd__nand4_1 _10609_ (.A(_05232_),
    .B(_05233_),
    .C(_05234_),
    .D(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__a22oi_1 _10610_ (.A1(\core.CPU_Dmem_value_a5[12][24] ),
    .A2(net524),
    .B1(net505),
    .B2(\core.CPU_Dmem_value_a5[3][24] ),
    .Y(_05237_));
 sky130_fd_sc_hd__a22oi_1 _10611_ (.A1(\core.CPU_Dmem_value_a5[2][24] ),
    .A2(net508),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][24] ),
    .Y(_05238_));
 sky130_fd_sc_hd__a22oi_1 _10612_ (.A1(\core.CPU_Dmem_value_a5[6][24] ),
    .A2(net492),
    .B1(_02428_),
    .B2(\core.CPU_Dmem_value_a5[9][24] ),
    .Y(_05239_));
 sky130_fd_sc_hd__a21oi_1 _10613_ (.A1(\core.CPU_Dmem_value_a5[8][24] ),
    .A2(net485),
    .B1(net558),
    .Y(_05240_));
 sky130_fd_sc_hd__nand4_1 _10614_ (.A(_05237_),
    .B(_05238_),
    .C(_05239_),
    .D(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__o22a_1 _10615_ (.A1(\core.CPU_Dmem_value_a5[0][24] ),
    .A2(net534),
    .B1(_05236_),
    .B2(_05241_),
    .X(\core.w_CPU_dmem_rd_data_a4[24] ));
 sky130_fd_sc_hd__a21oi_1 _10616_ (.A1(\core.CPU_Dmem_value_a5[4][25] ),
    .A2(net500),
    .B1(net559),
    .Y(_05242_));
 sky130_fd_sc_hd__a22oi_1 _10617_ (.A1(\core.CPU_Dmem_value_a5[11][25] ),
    .A2(net527),
    .B1(net518),
    .B2(\core.CPU_Dmem_value_a5[14][25] ),
    .Y(_05243_));
 sky130_fd_sc_hd__a22oi_1 _10618_ (.A1(\core.CPU_Dmem_value_a5[13][25] ),
    .A2(net522),
    .B1(net517),
    .B2(\core.CPU_Dmem_value_a5[15][25] ),
    .Y(_05244_));
 sky130_fd_sc_hd__a22oi_1 _10619_ (.A1(\core.CPU_Dmem_value_a5[10][25] ),
    .A2(net530),
    .B1(net523),
    .B2(\core.CPU_Dmem_value_a5[12][25] ),
    .Y(_05245_));
 sky130_fd_sc_hd__nand4_1 _10620_ (.A(_05242_),
    .B(_05243_),
    .C(_05244_),
    .D(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__a22o_1 _10621_ (.A1(\core.CPU_Dmem_value_a5[2][25] ),
    .A2(net508),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][25] ),
    .X(_05247_));
 sky130_fd_sc_hd__a221oi_1 _10622_ (.A1(\core.CPU_Dmem_value_a5[1][25] ),
    .A2(net514),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][25] ),
    .C1(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__a22oi_1 _10623_ (.A1(\core.CPU_Dmem_value_a5[3][25] ),
    .A2(net505),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][25] ),
    .Y(_05249_));
 sky130_fd_sc_hd__a22oi_1 _10624_ (.A1(\core.CPU_Dmem_value_a5[5][25] ),
    .A2(net497),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][25] ),
    .Y(_05250_));
 sky130_fd_sc_hd__nand3_1 _10625_ (.A(_05248_),
    .B(_05249_),
    .C(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__o22a_1 _10626_ (.A1(\core.CPU_Dmem_value_a5[0][25] ),
    .A2(net534),
    .B1(_05246_),
    .B2(_05251_),
    .X(\core.w_CPU_dmem_rd_data_a4[25] ));
 sky130_fd_sc_hd__a21oi_1 _10628_ (.A1(\core.CPU_Dmem_value_a5[5][26] ),
    .A2(net498),
    .B1(net559),
    .Y(_05253_));
 sky130_fd_sc_hd__a22oi_1 _10629_ (.A1(\core.CPU_Dmem_value_a5[12][26] ),
    .A2(net523),
    .B1(net514),
    .B2(\core.CPU_Dmem_value_a5[1][26] ),
    .Y(_05254_));
 sky130_fd_sc_hd__a22oi_1 _10630_ (.A1(\core.CPU_Dmem_value_a5[11][26] ),
    .A2(net528),
    .B1(net518),
    .B2(\core.CPU_Dmem_value_a5[14][26] ),
    .Y(_05255_));
 sky130_fd_sc_hd__a22oi_1 _10631_ (.A1(\core.CPU_Dmem_value_a5[10][26] ),
    .A2(net530),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][26] ),
    .Y(_05256_));
 sky130_fd_sc_hd__nand4_1 _10632_ (.A(_05253_),
    .B(_05254_),
    .C(_05255_),
    .D(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__a22o_1 _10633_ (.A1(\core.CPU_Dmem_value_a5[2][26] ),
    .A2(net508),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][26] ),
    .X(_05258_));
 sky130_fd_sc_hd__a221oi_1 _10634_ (.A1(\core.CPU_Dmem_value_a5[3][26] ),
    .A2(net506),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][26] ),
    .C1(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__a22oi_1 _10635_ (.A1(\core.CPU_Dmem_value_a5[13][26] ),
    .A2(net522),
    .B1(net484),
    .B2(\core.CPU_Dmem_value_a5[8][26] ),
    .Y(_05260_));
 sky130_fd_sc_hd__a22oi_1 _10636_ (.A1(\core.CPU_Dmem_value_a5[15][26] ),
    .A2(_01734_),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][26] ),
    .Y(_05261_));
 sky130_fd_sc_hd__nand3_1 _10637_ (.A(_05259_),
    .B(_05260_),
    .C(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__o22a_1 _10638_ (.A1(\core.CPU_Dmem_value_a5[0][26] ),
    .A2(net534),
    .B1(_05257_),
    .B2(_05262_),
    .X(\core.w_CPU_dmem_rd_data_a4[26] ));
 sky130_fd_sc_hd__a21oi_1 _10639_ (.A1(\core.CPU_Dmem_value_a5[8][27] ),
    .A2(net484),
    .B1(net559),
    .Y(_05263_));
 sky130_fd_sc_hd__a22oi_1 _10640_ (.A1(\core.CPU_Dmem_value_a5[12][27] ),
    .A2(net523),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][27] ),
    .Y(_05264_));
 sky130_fd_sc_hd__a22oi_1 _10641_ (.A1(\core.CPU_Dmem_value_a5[5][27] ),
    .A2(net498),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][27] ),
    .Y(_05265_));
 sky130_fd_sc_hd__a22oi_1 _10642_ (.A1(\core.CPU_Dmem_value_a5[14][27] ),
    .A2(_01660_),
    .B1(_01734_),
    .B2(\core.CPU_Dmem_value_a5[15][27] ),
    .Y(_05266_));
 sky130_fd_sc_hd__nand4_1 _10643_ (.A(_05263_),
    .B(_05264_),
    .C(_05265_),
    .D(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__a22o_1 _10644_ (.A1(\core.CPU_Dmem_value_a5[1][27] ),
    .A2(net514),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][27] ),
    .X(_05268_));
 sky130_fd_sc_hd__a221oi_1 _10645_ (.A1(\core.CPU_Dmem_value_a5[13][27] ),
    .A2(_01582_),
    .B1(net506),
    .B2(\core.CPU_Dmem_value_a5[3][27] ),
    .C1(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__a22oi_1 _10646_ (.A1(\core.CPU_Dmem_value_a5[10][27] ),
    .A2(net530),
    .B1(net507),
    .B2(\core.CPU_Dmem_value_a5[2][27] ),
    .Y(_05270_));
 sky130_fd_sc_hd__a22oi_1 _10647_ (.A1(\core.CPU_Dmem_value_a5[11][27] ),
    .A2(net528),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][27] ),
    .Y(_05271_));
 sky130_fd_sc_hd__nand3_1 _10648_ (.A(_05269_),
    .B(_05270_),
    .C(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__o22a_1 _10649_ (.A1(\core.CPU_Dmem_value_a5[0][27] ),
    .A2(_01199_),
    .B1(_05267_),
    .B2(_05272_),
    .X(\core.w_CPU_dmem_rd_data_a4[27] ));
 sky130_fd_sc_hd__a21oi_1 _10650_ (.A1(\core.CPU_Dmem_value_a5[2][28] ),
    .A2(net507),
    .B1(net559),
    .Y(_05273_));
 sky130_fd_sc_hd__a22oi_1 _10651_ (.A1(\core.CPU_Dmem_value_a5[10][28] ),
    .A2(net530),
    .B1(net517),
    .B2(\core.CPU_Dmem_value_a5[15][28] ),
    .Y(_05274_));
 sky130_fd_sc_hd__a22oi_1 _10652_ (.A1(\core.CPU_Dmem_value_a5[1][28] ),
    .A2(net514),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][28] ),
    .Y(_05275_));
 sky130_fd_sc_hd__a22oi_1 _10653_ (.A1(\core.CPU_Dmem_value_a5[12][28] ),
    .A2(net523),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][28] ),
    .Y(_05276_));
 sky130_fd_sc_hd__nand4_1 _10654_ (.A(_05273_),
    .B(_05274_),
    .C(_05275_),
    .D(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__a22oi_1 _10655_ (.A1(\core.CPU_Dmem_value_a5[11][28] ),
    .A2(net528),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][28] ),
    .Y(_05278_));
 sky130_fd_sc_hd__a22oi_1 _10656_ (.A1(\core.CPU_Dmem_value_a5[3][28] ),
    .A2(net506),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][28] ),
    .Y(_05279_));
 sky130_fd_sc_hd__a22oi_1 _10657_ (.A1(\core.CPU_Dmem_value_a5[14][28] ),
    .A2(net518),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][28] ),
    .Y(_05280_));
 sky130_fd_sc_hd__a22oi_1 _10658_ (.A1(\core.CPU_Dmem_value_a5[5][28] ),
    .A2(net498),
    .B1(net484),
    .B2(\core.CPU_Dmem_value_a5[8][28] ),
    .Y(_05281_));
 sky130_fd_sc_hd__nand4_1 _10659_ (.A(_05278_),
    .B(_05279_),
    .C(_05280_),
    .D(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__o22a_1 _10660_ (.A1(\core.CPU_Dmem_value_a5[0][28] ),
    .A2(net534),
    .B1(_05277_),
    .B2(_05282_),
    .X(\core.w_CPU_dmem_rd_data_a4[28] ));
 sky130_fd_sc_hd__a22oi_1 _10661_ (.A1(\core.CPU_Dmem_value_a5[12][29] ),
    .A2(net524),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][29] ),
    .Y(_05283_));
 sky130_fd_sc_hd__a22oi_1 _10662_ (.A1(\core.CPU_Dmem_value_a5[14][29] ),
    .A2(net518),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][29] ),
    .Y(_05284_));
 sky130_fd_sc_hd__a22oi_1 _10663_ (.A1(\core.CPU_Dmem_value_a5[1][29] ),
    .A2(net513),
    .B1(net497),
    .B2(\core.CPU_Dmem_value_a5[5][29] ),
    .Y(_05285_));
 sky130_fd_sc_hd__a22oi_1 _10664_ (.A1(\core.CPU_Dmem_value_a5[10][29] ),
    .A2(net529),
    .B1(_02275_),
    .B2(\core.CPU_Dmem_value_a5[7][29] ),
    .Y(_05286_));
 sky130_fd_sc_hd__nand4_1 _10665_ (.A(_05283_),
    .B(_05284_),
    .C(_05285_),
    .D(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__a22oi_1 _10666_ (.A1(\core.CPU_Dmem_value_a5[11][29] ),
    .A2(net527),
    .B1(net508),
    .B2(\core.CPU_Dmem_value_a5[2][29] ),
    .Y(_05288_));
 sky130_fd_sc_hd__a22oi_1 _10667_ (.A1(\core.CPU_Dmem_value_a5[3][29] ),
    .A2(net505),
    .B1(net499),
    .B2(\core.CPU_Dmem_value_a5[4][29] ),
    .Y(_05289_));
 sky130_fd_sc_hd__a22oi_1 _10668_ (.A1(\core.CPU_Dmem_value_a5[6][29] ),
    .A2(net491),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][29] ),
    .Y(_05290_));
 sky130_fd_sc_hd__a21oi_1 _10669_ (.A1(\core.CPU_Dmem_value_a5[15][29] ),
    .A2(net517),
    .B1(net558),
    .Y(_05291_));
 sky130_fd_sc_hd__nand4_1 _10670_ (.A(_05288_),
    .B(_05289_),
    .C(_05290_),
    .D(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__o22a_1 _10671_ (.A1(\core.CPU_Dmem_value_a5[0][29] ),
    .A2(net534),
    .B1(_05287_),
    .B2(_05292_),
    .X(\core.w_CPU_dmem_rd_data_a4[29] ));
 sky130_fd_sc_hd__a21oi_1 _10672_ (.A1(\core.CPU_Dmem_value_a5[8][2] ),
    .A2(net485),
    .B1(net559),
    .Y(_05293_));
 sky130_fd_sc_hd__a22oi_1 _10673_ (.A1(\core.CPU_Dmem_value_a5[13][2] ),
    .A2(net522),
    .B1(net518),
    .B2(\core.CPU_Dmem_value_a5[14][2] ),
    .Y(_05294_));
 sky130_fd_sc_hd__a22oi_1 _10674_ (.A1(\core.CPU_Dmem_value_a5[1][2] ),
    .A2(net514),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][2] ),
    .Y(_05295_));
 sky130_fd_sc_hd__a22oi_1 _10675_ (.A1(\core.CPU_Dmem_value_a5[11][2] ),
    .A2(net528),
    .B1(net517),
    .B2(\core.CPU_Dmem_value_a5[15][2] ),
    .Y(_05296_));
 sky130_fd_sc_hd__nand4_1 _10676_ (.A(_05293_),
    .B(_05294_),
    .C(_05295_),
    .D(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__a22oi_1 _10677_ (.A1(\core.CPU_Dmem_value_a5[10][2] ),
    .A2(net530),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][2] ),
    .Y(_05298_));
 sky130_fd_sc_hd__a22oi_1 _10678_ (.A1(\core.CPU_Dmem_value_a5[2][2] ),
    .A2(net507),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][2] ),
    .Y(_05299_));
 sky130_fd_sc_hd__a22oi_1 _10679_ (.A1(\core.CPU_Dmem_value_a5[12][2] ),
    .A2(net523),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][2] ),
    .Y(_05300_));
 sky130_fd_sc_hd__a22oi_1 _10680_ (.A1(\core.CPU_Dmem_value_a5[3][2] ),
    .A2(net506),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][2] ),
    .Y(_05301_));
 sky130_fd_sc_hd__nand4_1 _10681_ (.A(_05298_),
    .B(_05299_),
    .C(_05300_),
    .D(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__o22a_1 _10682_ (.A1(\core.CPU_Dmem_value_a5[0][2] ),
    .A2(net534),
    .B1(_05297_),
    .B2(_05302_),
    .X(\core.w_CPU_dmem_rd_data_a4[2] ));
 sky130_fd_sc_hd__a22oi_1 _10683_ (.A1(\core.CPU_Dmem_value_a5[14][30] ),
    .A2(net518),
    .B1(net517),
    .B2(\core.CPU_Dmem_value_a5[15][30] ),
    .Y(_05303_));
 sky130_fd_sc_hd__a22oi_1 _10684_ (.A1(\core.CPU_Dmem_value_a5[5][30] ),
    .A2(net497),
    .B1(net491),
    .B2(\core.CPU_Dmem_value_a5[6][30] ),
    .Y(_05304_));
 sky130_fd_sc_hd__a22oi_1 _10685_ (.A1(\core.CPU_Dmem_value_a5[10][30] ),
    .A2(net529),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][30] ),
    .Y(_05305_));
 sky130_fd_sc_hd__a22oi_1 _10686_ (.A1(\core.CPU_Dmem_value_a5[12][30] ),
    .A2(net524),
    .B1(_02275_),
    .B2(\core.CPU_Dmem_value_a5[7][30] ),
    .Y(_05306_));
 sky130_fd_sc_hd__nand4_1 _10687_ (.A(_05303_),
    .B(_05304_),
    .C(_05305_),
    .D(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__mux2i_1 _10688_ (.A0(\core.CPU_Dmem_value_a5[2][30] ),
    .A1(\core.CPU_Dmem_value_a5[3][30] ),
    .S(\core.CPU_dmem_addr_a4[0] ),
    .Y(_05308_));
 sky130_fd_sc_hd__o21ai_0 _10689_ (.A1(\core.CPU_Dmem_value_a5[1][30] ),
    .A2(_01580_),
    .B1(_01195_),
    .Y(_05309_));
 sky130_fd_sc_hd__a21oi_1 _10690_ (.A1(\core.CPU_dmem_addr_a4[1] ),
    .A2(_05308_),
    .B1(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__a22oi_1 _10691_ (.A1(\core.CPU_Dmem_value_a5[11][30] ),
    .A2(net527),
    .B1(net499),
    .B2(\core.CPU_Dmem_value_a5[4][30] ),
    .Y(_05311_));
 sky130_fd_sc_hd__a22oi_1 _10692_ (.A1(\core.CPU_Dmem_value_a5[13][30] ),
    .A2(net522),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][30] ),
    .Y(_05312_));
 sky130_fd_sc_hd__nand2_1 _10693_ (.A(_05311_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__o32a_1 _10694_ (.A1(_05307_),
    .A2(_05310_),
    .A3(_05313_),
    .B1(net534),
    .B2(\core.CPU_Dmem_value_a5[0][30] ),
    .X(\core.w_CPU_dmem_rd_data_a4[30] ));
 sky130_fd_sc_hd__a21oi_1 _10695_ (.A1(\core.CPU_Dmem_value_a5[1][31] ),
    .A2(net514),
    .B1(net558),
    .Y(_05314_));
 sky130_fd_sc_hd__a22oi_1 _10696_ (.A1(\core.CPU_Dmem_value_a5[12][31] ),
    .A2(net524),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][31] ),
    .Y(_05315_));
 sky130_fd_sc_hd__a22oi_1 _10697_ (.A1(\core.CPU_Dmem_value_a5[15][31] ),
    .A2(net517),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][31] ),
    .Y(_05316_));
 sky130_fd_sc_hd__a22oi_1 _10698_ (.A1(\core.CPU_Dmem_value_a5[10][31] ),
    .A2(net530),
    .B1(net518),
    .B2(\core.CPU_Dmem_value_a5[14][31] ),
    .Y(_05317_));
 sky130_fd_sc_hd__nand4_1 _10699_ (.A(_05314_),
    .B(_05315_),
    .C(_05316_),
    .D(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__a22oi_1 _10700_ (.A1(\core.CPU_Dmem_value_a5[11][31] ),
    .A2(net528),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][31] ),
    .Y(_05319_));
 sky130_fd_sc_hd__a22oi_1 _10701_ (.A1(\core.CPU_Dmem_value_a5[2][31] ),
    .A2(net508),
    .B1(net506),
    .B2(\core.CPU_Dmem_value_a5[3][31] ),
    .Y(_05320_));
 sky130_fd_sc_hd__a22oi_1 _10702_ (.A1(\core.CPU_Dmem_value_a5[6][31] ),
    .A2(net492),
    .B1(_02428_),
    .B2(\core.CPU_Dmem_value_a5[9][31] ),
    .Y(_05321_));
 sky130_fd_sc_hd__a22oi_1 _10703_ (.A1(\core.CPU_Dmem_value_a5[5][31] ),
    .A2(net498),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][31] ),
    .Y(_05322_));
 sky130_fd_sc_hd__nand4_1 _10704_ (.A(_05319_),
    .B(_05320_),
    .C(_05321_),
    .D(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__o22a_1 _10705_ (.A1(\core.CPU_Dmem_value_a5[0][31] ),
    .A2(net534),
    .B1(_05318_),
    .B2(_05323_),
    .X(\core.w_CPU_dmem_rd_data_a4[31] ));
 sky130_fd_sc_hd__a22o_1 _10706_ (.A1(\core.CPU_Dmem_value_a5[15][3] ),
    .A2(net517),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][3] ),
    .X(_05324_));
 sky130_fd_sc_hd__a221oi_1 _10707_ (.A1(\core.CPU_Dmem_value_a5[14][3] ),
    .A2(net518),
    .B1(net491),
    .B2(\core.CPU_Dmem_value_a5[6][3] ),
    .C1(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__a22oi_1 _10708_ (.A1(\core.CPU_Dmem_value_a5[11][3] ),
    .A2(net527),
    .B1(_02275_),
    .B2(\core.CPU_Dmem_value_a5[7][3] ),
    .Y(_05326_));
 sky130_fd_sc_hd__a22oi_1 _10709_ (.A1(\core.CPU_Dmem_value_a5[13][3] ),
    .A2(net522),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][3] ),
    .Y(_05327_));
 sky130_fd_sc_hd__and3_1 _10710_ (.A(_05325_),
    .B(_05326_),
    .C(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__mux2i_1 _10711_ (.A0(\core.CPU_Dmem_value_a5[2][3] ),
    .A1(\core.CPU_Dmem_value_a5[3][3] ),
    .S(\core.CPU_dmem_addr_a4[0] ),
    .Y(_05329_));
 sky130_fd_sc_hd__o21ai_0 _10712_ (.A1(\core.CPU_Dmem_value_a5[1][3] ),
    .A2(_01580_),
    .B1(_01195_),
    .Y(_05330_));
 sky130_fd_sc_hd__a21oi_1 _10713_ (.A1(\core.CPU_dmem_addr_a4[1] ),
    .A2(_05329_),
    .B1(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__a221oi_1 _10714_ (.A1(\core.CPU_Dmem_value_a5[10][3] ),
    .A2(net529),
    .B1(net499),
    .B2(\core.CPU_Dmem_value_a5[4][3] ),
    .C1(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__a22oi_1 _10715_ (.A1(\core.CPU_Dmem_value_a5[12][3] ),
    .A2(net523),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][3] ),
    .Y(_05333_));
 sky130_fd_sc_hd__nor2_1 _10716_ (.A(\core.CPU_Dmem_value_a5[0][3] ),
    .B(net534),
    .Y(_05334_));
 sky130_fd_sc_hd__a31oi_1 _10717_ (.A1(_05328_),
    .A2(_05332_),
    .A3(_05333_),
    .B1(_05334_),
    .Y(\core.w_CPU_dmem_rd_data_a4[3] ));
 sky130_fd_sc_hd__a21oi_1 _10718_ (.A1(\core.CPU_Dmem_value_a5[8][4] ),
    .A2(net484),
    .B1(net559),
    .Y(_05335_));
 sky130_fd_sc_hd__a22oi_1 _10719_ (.A1(\core.CPU_Dmem_value_a5[13][4] ),
    .A2(_01582_),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][4] ),
    .Y(_05336_));
 sky130_fd_sc_hd__a22oi_1 _10720_ (.A1(\core.CPU_Dmem_value_a5[12][4] ),
    .A2(net523),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][4] ),
    .Y(_05337_));
 sky130_fd_sc_hd__a22oi_1 _10721_ (.A1(\core.CPU_Dmem_value_a5[11][4] ),
    .A2(net528),
    .B1(net514),
    .B2(\core.CPU_Dmem_value_a5[1][4] ),
    .Y(_05338_));
 sky130_fd_sc_hd__nand4_1 _10722_ (.A(_05335_),
    .B(_05336_),
    .C(_05337_),
    .D(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__a22oi_1 _10723_ (.A1(\core.CPU_Dmem_value_a5[10][4] ),
    .A2(net529),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][4] ),
    .Y(_05340_));
 sky130_fd_sc_hd__a22oi_1 _10724_ (.A1(\core.CPU_Dmem_value_a5[15][4] ),
    .A2(_01734_),
    .B1(net507),
    .B2(\core.CPU_Dmem_value_a5[2][4] ),
    .Y(_05341_));
 sky130_fd_sc_hd__a22oi_1 _10725_ (.A1(\core.CPU_Dmem_value_a5[3][4] ),
    .A2(net506),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][4] ),
    .Y(_05342_));
 sky130_fd_sc_hd__a22oi_1 _10726_ (.A1(\core.CPU_Dmem_value_a5[14][4] ),
    .A2(_01660_),
    .B1(_02275_),
    .B2(\core.CPU_Dmem_value_a5[7][4] ),
    .Y(_05343_));
 sky130_fd_sc_hd__nand4_1 _10727_ (.A(_05340_),
    .B(_05341_),
    .C(_05342_),
    .D(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__o22a_1 _10728_ (.A1(\core.CPU_Dmem_value_a5[0][4] ),
    .A2(_01199_),
    .B1(_05339_),
    .B2(_05344_),
    .X(\core.w_CPU_dmem_rd_data_a4[4] ));
 sky130_fd_sc_hd__a21oi_1 _10729_ (.A1(\core.CPU_Dmem_value_a5[3][5] ),
    .A2(net506),
    .B1(net559),
    .Y(_05345_));
 sky130_fd_sc_hd__a22oi_1 _10730_ (.A1(\core.CPU_Dmem_value_a5[12][5] ),
    .A2(net523),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][5] ),
    .Y(_05346_));
 sky130_fd_sc_hd__a22oi_1 _10731_ (.A1(\core.CPU_Dmem_value_a5[13][5] ),
    .A2(_01582_),
    .B1(net484),
    .B2(\core.CPU_Dmem_value_a5[8][5] ),
    .Y(_05347_));
 sky130_fd_sc_hd__a22oi_1 _10732_ (.A1(\core.CPU_Dmem_value_a5[10][5] ),
    .A2(net530),
    .B1(_01734_),
    .B2(\core.CPU_Dmem_value_a5[15][5] ),
    .Y(_05348_));
 sky130_fd_sc_hd__nand4_1 _10733_ (.A(_05345_),
    .B(_05346_),
    .C(_05347_),
    .D(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__a22oi_1 _10734_ (.A1(\core.CPU_Dmem_value_a5[11][5] ),
    .A2(net528),
    .B1(net514),
    .B2(\core.CPU_Dmem_value_a5[1][5] ),
    .Y(_05350_));
 sky130_fd_sc_hd__a22oi_1 _10735_ (.A1(\core.CPU_Dmem_value_a5[2][5] ),
    .A2(net507),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][5] ),
    .Y(_05351_));
 sky130_fd_sc_hd__a22oi_1 _10736_ (.A1(\core.CPU_Dmem_value_a5[14][5] ),
    .A2(net518),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][5] ),
    .Y(_05352_));
 sky130_fd_sc_hd__a22oi_1 _10737_ (.A1(\core.CPU_Dmem_value_a5[5][5] ),
    .A2(net498),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][5] ),
    .Y(_05353_));
 sky130_fd_sc_hd__nand4_1 _10738_ (.A(_05350_),
    .B(_05351_),
    .C(_05352_),
    .D(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__o22a_1 _10739_ (.A1(\core.CPU_Dmem_value_a5[0][5] ),
    .A2(_01199_),
    .B1(_05349_),
    .B2(_05354_),
    .X(\core.w_CPU_dmem_rd_data_a4[5] ));
 sky130_fd_sc_hd__a21oi_1 _10740_ (.A1(\core.CPU_Dmem_value_a5[3][6] ),
    .A2(net505),
    .B1(net558),
    .Y(_05355_));
 sky130_fd_sc_hd__a22oi_1 _10741_ (.A1(\core.CPU_Dmem_value_a5[12][6] ),
    .A2(net524),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][6] ),
    .Y(_05356_));
 sky130_fd_sc_hd__a22oi_1 _10742_ (.A1(\core.CPU_Dmem_value_a5[15][6] ),
    .A2(net517),
    .B1(net513),
    .B2(\core.CPU_Dmem_value_a5[1][6] ),
    .Y(_05357_));
 sky130_fd_sc_hd__a22oi_1 _10743_ (.A1(\core.CPU_Dmem_value_a5[10][6] ),
    .A2(net529),
    .B1(net518),
    .B2(\core.CPU_Dmem_value_a5[14][6] ),
    .Y(_05358_));
 sky130_fd_sc_hd__nand4_1 _10744_ (.A(_05355_),
    .B(_05356_),
    .C(_05357_),
    .D(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__a22oi_1 _10745_ (.A1(\core.CPU_Dmem_value_a5[11][6] ),
    .A2(net527),
    .B1(net522),
    .B2(\core.CPU_Dmem_value_a5[13][6] ),
    .Y(_05360_));
 sky130_fd_sc_hd__a22oi_1 _10746_ (.A1(\core.CPU_Dmem_value_a5[2][6] ),
    .A2(net508),
    .B1(net499),
    .B2(\core.CPU_Dmem_value_a5[4][6] ),
    .Y(_05361_));
 sky130_fd_sc_hd__a22oi_1 _10747_ (.A1(\core.CPU_Dmem_value_a5[5][6] ),
    .A2(net497),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][6] ),
    .Y(_05362_));
 sky130_fd_sc_hd__a22oi_1 _10748_ (.A1(\core.CPU_Dmem_value_a5[6][6] ),
    .A2(net491),
    .B1(_02275_),
    .B2(\core.CPU_Dmem_value_a5[7][6] ),
    .Y(_05363_));
 sky130_fd_sc_hd__nand4_1 _10749_ (.A(_05360_),
    .B(_05361_),
    .C(_05362_),
    .D(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__o22a_1 _10750_ (.A1(\core.CPU_Dmem_value_a5[0][6] ),
    .A2(net534),
    .B1(_05359_),
    .B2(_05364_),
    .X(\core.w_CPU_dmem_rd_data_a4[6] ));
 sky130_fd_sc_hd__a21oi_1 _10751_ (.A1(\core.CPU_Dmem_value_a5[2][7] ),
    .A2(net508),
    .B1(net558),
    .Y(_05365_));
 sky130_fd_sc_hd__a22oi_1 _10752_ (.A1(\core.CPU_Dmem_value_a5[10][7] ),
    .A2(net529),
    .B1(net517),
    .B2(\core.CPU_Dmem_value_a5[15][7] ),
    .Y(_05366_));
 sky130_fd_sc_hd__a22oi_1 _10753_ (.A1(\core.CPU_Dmem_value_a5[1][7] ),
    .A2(net513),
    .B1(net497),
    .B2(\core.CPU_Dmem_value_a5[5][7] ),
    .Y(_05367_));
 sky130_fd_sc_hd__a22oi_1 _10754_ (.A1(\core.CPU_Dmem_value_a5[11][7] ),
    .A2(net527),
    .B1(net524),
    .B2(\core.CPU_Dmem_value_a5[12][7] ),
    .Y(_05368_));
 sky130_fd_sc_hd__nand4_1 _10755_ (.A(_05365_),
    .B(_05366_),
    .C(_05367_),
    .D(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__a22oi_1 _10756_ (.A1(\core.CPU_Dmem_value_a5[13][7] ),
    .A2(net522),
    .B1(net518),
    .B2(\core.CPU_Dmem_value_a5[14][7] ),
    .Y(_05370_));
 sky130_fd_sc_hd__a22oi_1 _10757_ (.A1(\core.CPU_Dmem_value_a5[3][7] ),
    .A2(net505),
    .B1(net499),
    .B2(\core.CPU_Dmem_value_a5[4][7] ),
    .Y(_05371_));
 sky130_fd_sc_hd__a22oi_1 _10758_ (.A1(\core.CPU_Dmem_value_a5[6][7] ),
    .A2(net491),
    .B1(net483),
    .B2(\core.CPU_Dmem_value_a5[9][7] ),
    .Y(_05372_));
 sky130_fd_sc_hd__a22oi_1 _10759_ (.A1(\core.CPU_Dmem_value_a5[7][7] ),
    .A2(_02275_),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][7] ),
    .Y(_05373_));
 sky130_fd_sc_hd__nand4_1 _10760_ (.A(_05370_),
    .B(_05371_),
    .C(_05372_),
    .D(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__o22a_1 _10761_ (.A1(\core.CPU_Dmem_value_a5[0][7] ),
    .A2(net534),
    .B1(_05369_),
    .B2(_05374_),
    .X(\core.w_CPU_dmem_rd_data_a4[7] ));
 sky130_fd_sc_hd__a21oi_1 _10762_ (.A1(\core.CPU_Dmem_value_a5[9][8] ),
    .A2(_02428_),
    .B1(net559),
    .Y(_05375_));
 sky130_fd_sc_hd__a22oi_1 _10763_ (.A1(\core.CPU_Dmem_value_a5[12][8] ),
    .A2(net524),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][8] ),
    .Y(_05376_));
 sky130_fd_sc_hd__a22oi_1 _10764_ (.A1(\core.CPU_Dmem_value_a5[11][8] ),
    .A2(net528),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][8] ),
    .Y(_05377_));
 sky130_fd_sc_hd__a22oi_1 _10765_ (.A1(\core.CPU_Dmem_value_a5[14][8] ),
    .A2(net518),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][8] ),
    .Y(_05378_));
 sky130_fd_sc_hd__nand4_1 _10766_ (.A(_05375_),
    .B(_05376_),
    .C(_05377_),
    .D(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__a22o_1 _10767_ (.A1(\core.CPU_Dmem_value_a5[2][8] ),
    .A2(net508),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][8] ),
    .X(_05380_));
 sky130_fd_sc_hd__a221oi_1 _10768_ (.A1(\core.CPU_Dmem_value_a5[15][8] ),
    .A2(net517),
    .B1(net505),
    .B2(\core.CPU_Dmem_value_a5[3][8] ),
    .C1(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__a22oi_1 _10769_ (.A1(\core.CPU_Dmem_value_a5[10][8] ),
    .A2(net530),
    .B1(net514),
    .B2(\core.CPU_Dmem_value_a5[1][8] ),
    .Y(_05382_));
 sky130_fd_sc_hd__a22oi_1 _10770_ (.A1(\core.CPU_Dmem_value_a5[13][8] ),
    .A2(net522),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][8] ),
    .Y(_05383_));
 sky130_fd_sc_hd__nand3_1 _10771_ (.A(_05381_),
    .B(_05382_),
    .C(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__o22a_1 _10772_ (.A1(\core.CPU_Dmem_value_a5[0][8] ),
    .A2(net534),
    .B1(_05379_),
    .B2(_05384_),
    .X(\core.w_CPU_dmem_rd_data_a4[8] ));
 sky130_fd_sc_hd__a21oi_1 _10773_ (.A1(\core.CPU_Dmem_value_a5[9][9] ),
    .A2(_02428_),
    .B1(net559),
    .Y(_05385_));
 sky130_fd_sc_hd__a22oi_1 _10774_ (.A1(\core.CPU_Dmem_value_a5[10][9] ),
    .A2(net530),
    .B1(net485),
    .B2(\core.CPU_Dmem_value_a5[8][9] ),
    .Y(_05386_));
 sky130_fd_sc_hd__a22oi_1 _10775_ (.A1(\core.CPU_Dmem_value_a5[12][9] ),
    .A2(net524),
    .B1(net498),
    .B2(\core.CPU_Dmem_value_a5[5][9] ),
    .Y(_05387_));
 sky130_fd_sc_hd__a22oi_1 _10776_ (.A1(\core.CPU_Dmem_value_a5[15][9] ),
    .A2(net517),
    .B1(net500),
    .B2(\core.CPU_Dmem_value_a5[4][9] ),
    .Y(_05388_));
 sky130_fd_sc_hd__nand4_1 _10777_ (.A(_05385_),
    .B(_05386_),
    .C(_05387_),
    .D(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__a22o_1 _10778_ (.A1(\core.CPU_Dmem_value_a5[3][9] ),
    .A2(net506),
    .B1(net490),
    .B2(\core.CPU_Dmem_value_a5[7][9] ),
    .X(_05390_));
 sky130_fd_sc_hd__a221oi_1 _10779_ (.A1(\core.CPU_Dmem_value_a5[14][9] ),
    .A2(net518),
    .B1(net514),
    .B2(\core.CPU_Dmem_value_a5[1][9] ),
    .C1(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__a22oi_1 _10780_ (.A1(\core.CPU_Dmem_value_a5[11][9] ),
    .A2(net528),
    .B1(net507),
    .B2(\core.CPU_Dmem_value_a5[2][9] ),
    .Y(_05392_));
 sky130_fd_sc_hd__a22oi_1 _10781_ (.A1(\core.CPU_Dmem_value_a5[13][9] ),
    .A2(net522),
    .B1(net492),
    .B2(\core.CPU_Dmem_value_a5[6][9] ),
    .Y(_05393_));
 sky130_fd_sc_hd__nand3_1 _10782_ (.A(_05391_),
    .B(_05392_),
    .C(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__o22a_1 _10783_ (.A1(\core.CPU_Dmem_value_a5[0][9] ),
    .A2(net534),
    .B1(_05389_),
    .B2(_05394_),
    .X(\core.w_CPU_dmem_rd_data_a4[9] ));
 sky130_fd_sc_hd__fa_1 _10784_ (.A(\core.CPU_imm_a3[1] ),
    .B(\core.CPU_src1_value_a3[1] ),
    .CIN(_00000_),
    .COUT(_00001_),
    .SUM(_00002_));
 sky130_fd_sc_hd__fa_1 _10785_ (.A(_00003_),
    .B(\core.CPU_src2_value_a3[1] ),
    .CIN(_00004_),
    .COUT(_00005_),
    .SUM(_00006_));
 sky130_fd_sc_hd__fa_1 _10786_ (.A(\core.CPU_src1_value_a3[1] ),
    .B(\core.CPU_src2_value_a3[1] ),
    .CIN(_00007_),
    .COUT(_00008_),
    .SUM(_00009_));
 sky130_fd_sc_hd__fa_1 _10787_ (.A(_00010_),
    .B(_00011_),
    .CIN(_00012_),
    .COUT(_00013_),
    .SUM(_00014_));
 sky130_fd_sc_hd__ha_1 _10788_ (.A(\core.CPU_imm_a2[1] ),
    .B(\core.CPU_inc_pc_a2[1] ),
    .COUT(_00015_),
    .SUM(_00016_));
 sky130_fd_sc_hd__ha_1 _10789_ (.A(\core.CPU_imm_a2[3] ),
    .B(\core.CPU_pc_a2[3] ),
    .COUT(_00017_),
    .SUM(_00018_));
 sky130_fd_sc_hd__ha_1 _10790_ (.A(\core.CPU_imm_a2[4] ),
    .B(\core.CPU_pc_a2[4] ),
    .COUT(_00019_),
    .SUM(_00020_));
 sky130_fd_sc_hd__ha_1 _10791_ (.A(_00021_),
    .B(\core.CPU_src2_value_a3[0] ),
    .COUT(_00004_),
    .SUM(_00022_));
 sky130_fd_sc_hd__ha_1 _10792_ (.A(\core.CPU_src1_value_a3[0] ),
    .B(\core.CPU_src2_value_a3[0] ),
    .COUT(_00007_),
    .SUM(_05395_));
 sky130_fd_sc_hd__ha_1 _10793_ (.A(\core.CPU_src1_value_a3[28] ),
    .B(_00023_),
    .COUT(_00024_),
    .SUM(_00025_));
 sky130_fd_sc_hd__ha_1 _10794_ (.A(\core.CPU_src1_value_a3[28] ),
    .B(\core.CPU_src2_value_a3[28] ),
    .COUT(_00026_),
    .SUM(_05396_));
 sky130_fd_sc_hd__ha_1 _10795_ (.A(\core.CPU_src1_value_a3[27] ),
    .B(_00027_),
    .COUT(_00028_),
    .SUM(_00029_));
 sky130_fd_sc_hd__ha_1 _10796_ (.A(\core.CPU_src1_value_a3[27] ),
    .B(\core.CPU_src2_value_a3[27] ),
    .COUT(_00030_),
    .SUM(_05397_));
 sky130_fd_sc_hd__ha_1 _10797_ (.A(\core.CPU_imm_a3[0] ),
    .B(\core.CPU_src1_value_a3[0] ),
    .COUT(_00000_),
    .SUM(_00031_));
 sky130_fd_sc_hd__ha_1 _10798_ (.A(\core.CPU_imm_a3[1] ),
    .B(\core.CPU_src1_value_a3[1] ),
    .COUT(_00032_),
    .SUM(_00033_));
 sky130_fd_sc_hd__ha_1 _10799_ (.A(\core.CPU_src1_value_a3[1] ),
    .B(_00035_),
    .COUT(_00036_),
    .SUM(_00034_));
 sky130_fd_sc_hd__ha_1 _10800_ (.A(\core.CPU_src1_value_a3[1] ),
    .B(\core.CPU_src2_value_a3[1] ),
    .COUT(_00037_),
    .SUM(_05398_));
 sky130_fd_sc_hd__ha_1 _10801_ (.A(\core.CPU_src1_value_a3[2] ),
    .B(_00038_),
    .COUT(_00039_),
    .SUM(_00040_));
 sky130_fd_sc_hd__ha_1 _10802_ (.A(\core.CPU_src1_value_a3[2] ),
    .B(\core.CPU_src2_value_a3[2] ),
    .COUT(_00041_),
    .SUM(_05399_));
 sky130_fd_sc_hd__ha_1 _10803_ (.A(\core.CPU_imm_a3[3] ),
    .B(\core.CPU_src1_value_a3[3] ),
    .COUT(_00042_),
    .SUM(_00043_));
 sky130_fd_sc_hd__ha_1 _10804_ (.A(\core.CPU_src1_value_a3[3] ),
    .B(_00044_),
    .COUT(_00045_),
    .SUM(_00046_));
 sky130_fd_sc_hd__ha_1 _10805_ (.A(\core.CPU_src1_value_a3[3] ),
    .B(\core.CPU_src2_value_a3[3] ),
    .COUT(_00047_),
    .SUM(_05400_));
 sky130_fd_sc_hd__ha_1 _10806_ (.A(\core.CPU_imm_a3[4] ),
    .B(\core.CPU_src1_value_a3[4] ),
    .COUT(_00048_),
    .SUM(_00049_));
 sky130_fd_sc_hd__ha_1 _10807_ (.A(\core.CPU_src1_value_a3[4] ),
    .B(_00050_),
    .COUT(_00051_),
    .SUM(_00052_));
 sky130_fd_sc_hd__ha_1 _10808_ (.A(\core.CPU_src1_value_a3[4] ),
    .B(\core.CPU_src2_value_a3[4] ),
    .COUT(_00053_),
    .SUM(_05401_));
 sky130_fd_sc_hd__ha_1 _10809_ (.A(\core.CPU_src1_value_a3[5] ),
    .B(_00054_),
    .COUT(_00055_),
    .SUM(_00056_));
 sky130_fd_sc_hd__ha_1 _10810_ (.A(\core.CPU_src1_value_a3[5] ),
    .B(\core.CPU_src2_value_a3[5] ),
    .COUT(_00057_),
    .SUM(_05402_));
 sky130_fd_sc_hd__ha_1 _10811_ (.A(\core.CPU_imm_a3[5] ),
    .B(\core.CPU_src1_value_a3[5] ),
    .COUT(_00058_),
    .SUM(_00059_));
 sky130_fd_sc_hd__ha_1 _10812_ (.A(\core.CPU_src1_value_a3[6] ),
    .B(_00060_),
    .COUT(_00061_),
    .SUM(_00062_));
 sky130_fd_sc_hd__ha_1 _10813_ (.A(\core.CPU_src1_value_a3[6] ),
    .B(\core.CPU_src2_value_a3[6] ),
    .COUT(_00063_),
    .SUM(_05403_));
 sky130_fd_sc_hd__ha_1 _10814_ (.A(net613),
    .B(\core.CPU_src1_value_a3[7] ),
    .COUT(_00064_),
    .SUM(_00065_));
 sky130_fd_sc_hd__ha_1 _10815_ (.A(net613),
    .B(\core.CPU_src1_value_a3[6] ),
    .COUT(_00066_),
    .SUM(_00067_));
 sky130_fd_sc_hd__ha_1 _10816_ (.A(\core.CPU_src1_value_a3[7] ),
    .B(_00068_),
    .COUT(_00069_),
    .SUM(_00070_));
 sky130_fd_sc_hd__ha_1 _10817_ (.A(\core.CPU_src1_value_a3[7] ),
    .B(\core.CPU_src2_value_a3[7] ),
    .COUT(_00071_),
    .SUM(_05404_));
 sky130_fd_sc_hd__ha_1 _10818_ (.A(net613),
    .B(\core.CPU_src1_value_a3[8] ),
    .COUT(_00072_),
    .SUM(_00073_));
 sky130_fd_sc_hd__ha_1 _10819_ (.A(\core.CPU_src1_value_a3[8] ),
    .B(_00074_),
    .COUT(_00075_),
    .SUM(_00076_));
 sky130_fd_sc_hd__ha_1 _10820_ (.A(\core.CPU_src1_value_a3[8] ),
    .B(\core.CPU_src2_value_a3[8] ),
    .COUT(_00077_),
    .SUM(_05405_));
 sky130_fd_sc_hd__ha_1 _10821_ (.A(\core.CPU_src1_value_a3[9] ),
    .B(_00078_),
    .COUT(_00079_),
    .SUM(_00080_));
 sky130_fd_sc_hd__ha_1 _10822_ (.A(\core.CPU_src1_value_a3[9] ),
    .B(\core.CPU_src2_value_a3[9] ),
    .COUT(_00081_),
    .SUM(_05406_));
 sky130_fd_sc_hd__ha_1 _10823_ (.A(net613),
    .B(\core.CPU_src1_value_a3[9] ),
    .COUT(_00082_),
    .SUM(_00083_));
 sky130_fd_sc_hd__ha_1 _10824_ (.A(\core.CPU_src1_value_a3[10] ),
    .B(_00084_),
    .COUT(_00085_),
    .SUM(_00086_));
 sky130_fd_sc_hd__ha_1 _10825_ (.A(\core.CPU_src1_value_a3[10] ),
    .B(\core.CPU_src2_value_a3[10] ),
    .COUT(_00087_),
    .SUM(_05407_));
 sky130_fd_sc_hd__ha_1 _10826_ (.A(\core.CPU_imm_a3[10] ),
    .B(\core.CPU_src1_value_a3[10] ),
    .COUT(_00088_),
    .SUM(_00089_));
 sky130_fd_sc_hd__ha_1 _10827_ (.A(\core.CPU_src1_value_a3[11] ),
    .B(_00090_),
    .COUT(_00091_),
    .SUM(_00092_));
 sky130_fd_sc_hd__ha_1 _10828_ (.A(\core.CPU_src1_value_a3[11] ),
    .B(\core.CPU_src2_value_a3[11] ),
    .COUT(_00093_),
    .SUM(_05408_));
 sky130_fd_sc_hd__ha_1 _10829_ (.A(\core.CPU_imm_a3[11] ),
    .B(\core.CPU_src1_value_a3[11] ),
    .COUT(_00094_),
    .SUM(_00095_));
 sky130_fd_sc_hd__ha_1 _10830_ (.A(\core.CPU_src1_value_a3[12] ),
    .B(_00096_),
    .COUT(_00097_),
    .SUM(_00098_));
 sky130_fd_sc_hd__ha_1 _10831_ (.A(\core.CPU_src1_value_a3[12] ),
    .B(\core.CPU_src2_value_a3[12] ),
    .COUT(_00099_),
    .SUM(_05409_));
 sky130_fd_sc_hd__ha_1 _10832_ (.A(net613),
    .B(\core.CPU_src1_value_a3[12] ),
    .COUT(_00100_),
    .SUM(_00101_));
 sky130_fd_sc_hd__ha_1 _10833_ (.A(\core.CPU_src1_value_a3[13] ),
    .B(_00102_),
    .COUT(_00103_),
    .SUM(_00104_));
 sky130_fd_sc_hd__ha_1 _10834_ (.A(\core.CPU_src1_value_a3[13] ),
    .B(\core.CPU_src2_value_a3[13] ),
    .COUT(_00105_),
    .SUM(_05410_));
 sky130_fd_sc_hd__ha_1 _10835_ (.A(net613),
    .B(\core.CPU_src1_value_a3[13] ),
    .COUT(_00106_),
    .SUM(_00107_));
 sky130_fd_sc_hd__ha_1 _10836_ (.A(\core.CPU_src1_value_a3[14] ),
    .B(_00108_),
    .COUT(_00109_),
    .SUM(_00110_));
 sky130_fd_sc_hd__ha_1 _10837_ (.A(\core.CPU_src1_value_a3[14] ),
    .B(\core.CPU_src2_value_a3[14] ),
    .COUT(_00111_),
    .SUM(_05411_));
 sky130_fd_sc_hd__ha_1 _10838_ (.A(net613),
    .B(\core.CPU_src1_value_a3[14] ),
    .COUT(_00112_),
    .SUM(_00113_));
 sky130_fd_sc_hd__ha_1 _10839_ (.A(\core.CPU_src1_value_a3[15] ),
    .B(_00114_),
    .COUT(_00115_),
    .SUM(_00116_));
 sky130_fd_sc_hd__ha_1 _10840_ (.A(\core.CPU_src1_value_a3[15] ),
    .B(\core.CPU_src2_value_a3[15] ),
    .COUT(_00117_),
    .SUM(_05412_));
 sky130_fd_sc_hd__ha_1 _10841_ (.A(net613),
    .B(\core.CPU_src1_value_a3[16] ),
    .COUT(_00118_),
    .SUM(_00119_));
 sky130_fd_sc_hd__ha_1 _10842_ (.A(net613),
    .B(\core.CPU_src1_value_a3[15] ),
    .COUT(_00120_),
    .SUM(_00121_));
 sky130_fd_sc_hd__ha_1 _10843_ (.A(\core.CPU_src1_value_a3[16] ),
    .B(_00122_),
    .COUT(_00123_),
    .SUM(_00124_));
 sky130_fd_sc_hd__ha_1 _10844_ (.A(\core.CPU_src1_value_a3[16] ),
    .B(\core.CPU_src2_value_a3[16] ),
    .COUT(_00125_),
    .SUM(_05413_));
 sky130_fd_sc_hd__ha_1 _10845_ (.A(net613),
    .B(\core.CPU_src1_value_a3[17] ),
    .COUT(_00126_),
    .SUM(_00127_));
 sky130_fd_sc_hd__ha_1 _10846_ (.A(\core.CPU_src1_value_a3[17] ),
    .B(_00128_),
    .COUT(_00129_),
    .SUM(_00130_));
 sky130_fd_sc_hd__ha_1 _10847_ (.A(\core.CPU_src1_value_a3[17] ),
    .B(\core.CPU_src2_value_a3[17] ),
    .COUT(_00131_),
    .SUM(_05414_));
 sky130_fd_sc_hd__ha_1 _10848_ (.A(net613),
    .B(\core.CPU_src1_value_a3[18] ),
    .COUT(_00132_),
    .SUM(_00133_));
 sky130_fd_sc_hd__ha_1 _10849_ (.A(\core.CPU_src1_value_a3[18] ),
    .B(_00134_),
    .COUT(_00135_),
    .SUM(_00136_));
 sky130_fd_sc_hd__ha_1 _10850_ (.A(\core.CPU_src1_value_a3[18] ),
    .B(\core.CPU_src2_value_a3[18] ),
    .COUT(_00137_),
    .SUM(_05415_));
 sky130_fd_sc_hd__ha_1 _10851_ (.A(net613),
    .B(\core.CPU_src1_value_a3[19] ),
    .COUT(_00138_),
    .SUM(_00139_));
 sky130_fd_sc_hd__ha_1 _10852_ (.A(\core.CPU_src1_value_a3[19] ),
    .B(_00140_),
    .COUT(_00141_),
    .SUM(_00142_));
 sky130_fd_sc_hd__ha_1 _10853_ (.A(\core.CPU_src1_value_a3[19] ),
    .B(\core.CPU_src2_value_a3[19] ),
    .COUT(_00143_),
    .SUM(_05416_));
 sky130_fd_sc_hd__ha_1 _10854_ (.A(net613),
    .B(\core.CPU_src1_value_a3[20] ),
    .COUT(_00144_),
    .SUM(_00145_));
 sky130_fd_sc_hd__ha_1 _10855_ (.A(\core.CPU_src1_value_a3[20] ),
    .B(_00146_),
    .COUT(_00147_),
    .SUM(_00148_));
 sky130_fd_sc_hd__ha_1 _10856_ (.A(\core.CPU_src1_value_a3[20] ),
    .B(\core.CPU_src2_value_a3[20] ),
    .COUT(_00149_),
    .SUM(_05417_));
 sky130_fd_sc_hd__ha_1 _10857_ (.A(net613),
    .B(\core.CPU_src1_value_a3[21] ),
    .COUT(_00150_),
    .SUM(_00151_));
 sky130_fd_sc_hd__ha_1 _10858_ (.A(\core.CPU_src1_value_a3[21] ),
    .B(_00152_),
    .COUT(_00153_),
    .SUM(_00154_));
 sky130_fd_sc_hd__ha_1 _10859_ (.A(\core.CPU_src1_value_a3[21] ),
    .B(\core.CPU_src2_value_a3[21] ),
    .COUT(_00155_),
    .SUM(_05418_));
 sky130_fd_sc_hd__ha_1 _10860_ (.A(net613),
    .B(\core.CPU_src1_value_a3[22] ),
    .COUT(_00156_),
    .SUM(_00157_));
 sky130_fd_sc_hd__ha_1 _10861_ (.A(\core.CPU_src1_value_a3[22] ),
    .B(_00158_),
    .COUT(_00159_),
    .SUM(_00160_));
 sky130_fd_sc_hd__ha_1 _10862_ (.A(\core.CPU_src1_value_a3[22] ),
    .B(\core.CPU_src2_value_a3[22] ),
    .COUT(_00161_),
    .SUM(_05419_));
 sky130_fd_sc_hd__ha_1 _10863_ (.A(net613),
    .B(\core.CPU_src1_value_a3[23] ),
    .COUT(_00162_),
    .SUM(_00163_));
 sky130_fd_sc_hd__ha_1 _10864_ (.A(\core.CPU_src1_value_a3[23] ),
    .B(_00164_),
    .COUT(_00165_),
    .SUM(_00166_));
 sky130_fd_sc_hd__ha_1 _10865_ (.A(\core.CPU_src1_value_a3[23] ),
    .B(\core.CPU_src2_value_a3[23] ),
    .COUT(_00167_),
    .SUM(_05420_));
 sky130_fd_sc_hd__ha_1 _10866_ (.A(net613),
    .B(\core.CPU_src1_value_a3[24] ),
    .COUT(_00168_),
    .SUM(_00169_));
 sky130_fd_sc_hd__ha_1 _10867_ (.A(\core.CPU_src1_value_a3[24] ),
    .B(_00170_),
    .COUT(_00171_),
    .SUM(_00172_));
 sky130_fd_sc_hd__ha_1 _10868_ (.A(\core.CPU_src1_value_a3[24] ),
    .B(\core.CPU_src2_value_a3[24] ),
    .COUT(_00173_),
    .SUM(_05421_));
 sky130_fd_sc_hd__ha_1 _10869_ (.A(net613),
    .B(\core.CPU_src1_value_a3[25] ),
    .COUT(_00174_),
    .SUM(_00175_));
 sky130_fd_sc_hd__ha_1 _10870_ (.A(\core.CPU_src1_value_a3[25] ),
    .B(_00176_),
    .COUT(_00177_),
    .SUM(_00178_));
 sky130_fd_sc_hd__ha_1 _10871_ (.A(\core.CPU_src1_value_a3[25] ),
    .B(\core.CPU_src2_value_a3[25] ),
    .COUT(_00179_),
    .SUM(_05422_));
 sky130_fd_sc_hd__ha_1 _10872_ (.A(net613),
    .B(\core.CPU_src1_value_a3[26] ),
    .COUT(_00180_),
    .SUM(_00181_));
 sky130_fd_sc_hd__ha_1 _10873_ (.A(\core.CPU_src1_value_a3[26] ),
    .B(_00182_),
    .COUT(_00183_),
    .SUM(_00184_));
 sky130_fd_sc_hd__ha_1 _10874_ (.A(\core.CPU_src1_value_a3[26] ),
    .B(\core.CPU_src2_value_a3[26] ),
    .COUT(_00185_),
    .SUM(_05423_));
 sky130_fd_sc_hd__ha_1 _10875_ (.A(net613),
    .B(\core.CPU_src1_value_a3[27] ),
    .COUT(_00186_),
    .SUM(_00187_));
 sky130_fd_sc_hd__ha_1 _10876_ (.A(net613),
    .B(\core.CPU_src1_value_a3[28] ),
    .COUT(_00188_),
    .SUM(_00189_));
 sky130_fd_sc_hd__ha_1 _10877_ (.A(net613),
    .B(\core.CPU_src1_value_a3[29] ),
    .COUT(_00190_),
    .SUM(_00191_));
 sky130_fd_sc_hd__ha_1 _10878_ (.A(\core.CPU_src1_value_a3[29] ),
    .B(_00192_),
    .COUT(_00193_),
    .SUM(_00194_));
 sky130_fd_sc_hd__ha_1 _10879_ (.A(\core.CPU_src1_value_a3[29] ),
    .B(net586),
    .COUT(_00195_),
    .SUM(_05424_));
 sky130_fd_sc_hd__ha_1 _10880_ (.A(net613),
    .B(\core.CPU_src1_value_a3[30] ),
    .COUT(_00196_),
    .SUM(_00197_));
 sky130_fd_sc_hd__ha_1 _10881_ (.A(\core.CPU_src1_value_a3[30] ),
    .B(_00198_),
    .COUT(_00199_),
    .SUM(_00200_));
 sky130_fd_sc_hd__ha_1 _10882_ (.A(\core.CPU_src1_value_a3[30] ),
    .B(\core.CPU_src2_value_a3[30] ),
    .COUT(_00201_),
    .SUM(_05425_));
 sky130_fd_sc_hd__ha_1 _10883_ (.A(\core.CPU_imm_a2[0] ),
    .B(\core.CPU_inc_pc_a2[0] ),
    .COUT(_00202_),
    .SUM(\core.CPU_br_tgt_pc_a2[0] ));
 sky130_fd_sc_hd__ha_1 _10884_ (.A(\core.CPU_inc_pc_a1[2] ),
    .B(_00203_),
    .COUT(_00204_),
    .SUM(\core.CPU_inc_pc_a1[3] ));
 sky130_fd_sc_hd__ha_1 _10885_ (.A(\core.CPU_inc_pc_a1[2] ),
    .B(\core.CPU_imem_rd_addr_a1[1] ),
    .COUT(_00205_),
    .SUM(_05426_));
 sky130_fd_sc_hd__ha_1 _10886_ (.A(\core.CPU_imem_rd_addr_a1[0] ),
    .B(_00203_),
    .COUT(_00206_),
    .SUM(_05427_));
 sky130_fd_sc_hd__ha_1 _10887_ (.A(\core.CPU_imem_rd_addr_a1[0] ),
    .B(\core.CPU_imem_rd_addr_a1[1] ),
    .COUT(_00207_),
    .SUM(_05428_));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][0]$_SDFFE_PP0P_  (.D(_00208_),
    .Q(\core.CPU_Dmem_value_a5[0][0] ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][10]$_SDFFE_PP0P_  (.D(_00209_),
    .Q(\core.CPU_Dmem_value_a5[0][10] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][11]$_SDFFE_PP0P_  (.D(_00210_),
    .Q(\core.CPU_Dmem_value_a5[0][11] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][12]$_SDFFE_PP0P_  (.D(_00211_),
    .Q(\core.CPU_Dmem_value_a5[0][12] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][13]$_SDFFE_PP0P_  (.D(_00212_),
    .Q(\core.CPU_Dmem_value_a5[0][13] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][14]$_SDFFE_PP0P_  (.D(_00213_),
    .Q(\core.CPU_Dmem_value_a5[0][14] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][15]$_SDFFE_PP0P_  (.D(_00214_),
    .Q(\core.CPU_Dmem_value_a5[0][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][16]$_SDFFE_PP0P_  (.D(_00215_),
    .Q(\core.CPU_Dmem_value_a5[0][16] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][17]$_SDFFE_PP0P_  (.D(_00216_),
    .Q(\core.CPU_Dmem_value_a5[0][17] ),
    .CLK(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][18]$_SDFFE_PP0P_  (.D(_00217_),
    .Q(\core.CPU_Dmem_value_a5[0][18] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][19]$_SDFFE_PP0P_  (.D(_00218_),
    .Q(\core.CPU_Dmem_value_a5[0][19] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][1]$_SDFFE_PP0P_  (.D(_00219_),
    .Q(\core.CPU_Dmem_value_a5[0][1] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][20]$_SDFFE_PP0P_  (.D(_00220_),
    .Q(\core.CPU_Dmem_value_a5[0][20] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][21]$_SDFFE_PP0P_  (.D(_00221_),
    .Q(\core.CPU_Dmem_value_a5[0][21] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][22]$_SDFFE_PP0P_  (.D(_00222_),
    .Q(\core.CPU_Dmem_value_a5[0][22] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][23]$_SDFFE_PP0P_  (.D(_00223_),
    .Q(\core.CPU_Dmem_value_a5[0][23] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][24]$_SDFFE_PP0P_  (.D(_00224_),
    .Q(\core.CPU_Dmem_value_a5[0][24] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][25]$_SDFFE_PP0P_  (.D(_00225_),
    .Q(\core.CPU_Dmem_value_a5[0][25] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][26]$_SDFFE_PP0P_  (.D(_00226_),
    .Q(\core.CPU_Dmem_value_a5[0][26] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][27]$_SDFFE_PP0P_  (.D(_00227_),
    .Q(\core.CPU_Dmem_value_a5[0][27] ),
    .CLK(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][28]$_SDFFE_PP0P_  (.D(_00228_),
    .Q(\core.CPU_Dmem_value_a5[0][28] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][29]$_SDFFE_PP0P_  (.D(_00229_),
    .Q(\core.CPU_Dmem_value_a5[0][29] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][2]$_SDFFE_PP0P_  (.D(_00230_),
    .Q(\core.CPU_Dmem_value_a5[0][2] ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][30]$_SDFFE_PP0P_  (.D(_00231_),
    .Q(\core.CPU_Dmem_value_a5[0][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][31]$_SDFFE_PP0P_  (.D(_00232_),
    .Q(\core.CPU_Dmem_value_a5[0][31] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][3]$_SDFFE_PP0P_  (.D(_00233_),
    .Q(\core.CPU_Dmem_value_a5[0][3] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][4]$_SDFFE_PP0P_  (.D(_00234_),
    .Q(\core.CPU_Dmem_value_a5[0][4] ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][5]$_SDFFE_PP0P_  (.D(_00235_),
    .Q(\core.CPU_Dmem_value_a5[0][5] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][6]$_SDFFE_PP0P_  (.D(_00236_),
    .Q(\core.CPU_Dmem_value_a5[0][6] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][7]$_SDFFE_PP0P_  (.D(_00237_),
    .Q(\core.CPU_Dmem_value_a5[0][7] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][8]$_SDFFE_PP0P_  (.D(_00238_),
    .Q(\core.CPU_Dmem_value_a5[0][8] ),
    .CLK(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[0][9]$_SDFFE_PP0P_  (.D(_00239_),
    .Q(\core.CPU_Dmem_value_a5[0][9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][0]$_SDFFE_PP0P_  (.D(_00240_),
    .Q(\core.CPU_Dmem_value_a5[10][0] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][10]$_SDFFE_PP0P_  (.D(_00241_),
    .Q(\core.CPU_Dmem_value_a5[10][10] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][11]$_SDFFE_PP0P_  (.D(_00242_),
    .Q(\core.CPU_Dmem_value_a5[10][11] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][12]$_SDFFE_PP0P_  (.D(_00243_),
    .Q(\core.CPU_Dmem_value_a5[10][12] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][13]$_SDFFE_PP0P_  (.D(_00244_),
    .Q(\core.CPU_Dmem_value_a5[10][13] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][14]$_SDFFE_PP0P_  (.D(_00245_),
    .Q(\core.CPU_Dmem_value_a5[10][14] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][15]$_SDFFE_PP0P_  (.D(_00246_),
    .Q(\core.CPU_Dmem_value_a5[10][15] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][16]$_SDFFE_PP0P_  (.D(_00247_),
    .Q(\core.CPU_Dmem_value_a5[10][16] ),
    .CLK(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][17]$_SDFFE_PP0P_  (.D(_00248_),
    .Q(\core.CPU_Dmem_value_a5[10][17] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][18]$_SDFFE_PP0P_  (.D(_00249_),
    .Q(\core.CPU_Dmem_value_a5[10][18] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][19]$_SDFFE_PP0P_  (.D(_00250_),
    .Q(\core.CPU_Dmem_value_a5[10][19] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][1]$_SDFFE_PP1P_  (.D(_00251_),
    .Q(\core.CPU_Dmem_value_a5[10][1] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][20]$_SDFFE_PP0P_  (.D(_00252_),
    .Q(\core.CPU_Dmem_value_a5[10][20] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][21]$_SDFFE_PP0P_  (.D(_00253_),
    .Q(\core.CPU_Dmem_value_a5[10][21] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][22]$_SDFFE_PP0P_  (.D(_00254_),
    .Q(\core.CPU_Dmem_value_a5[10][22] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][23]$_SDFFE_PP0P_  (.D(_00255_),
    .Q(\core.CPU_Dmem_value_a5[10][23] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][24]$_SDFFE_PP0P_  (.D(_00256_),
    .Q(\core.CPU_Dmem_value_a5[10][24] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][25]$_SDFFE_PP0P_  (.D(_00257_),
    .Q(\core.CPU_Dmem_value_a5[10][25] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][26]$_SDFFE_PP0P_  (.D(_00258_),
    .Q(\core.CPU_Dmem_value_a5[10][26] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][27]$_SDFFE_PP0P_  (.D(_00259_),
    .Q(\core.CPU_Dmem_value_a5[10][27] ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][28]$_SDFFE_PP0P_  (.D(_00260_),
    .Q(\core.CPU_Dmem_value_a5[10][28] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][29]$_SDFFE_PP0P_  (.D(_00261_),
    .Q(\core.CPU_Dmem_value_a5[10][29] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][2]$_SDFFE_PP0P_  (.D(_00262_),
    .Q(\core.CPU_Dmem_value_a5[10][2] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][30]$_SDFFE_PP0P_  (.D(_00263_),
    .Q(\core.CPU_Dmem_value_a5[10][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][31]$_SDFFE_PP0P_  (.D(_00264_),
    .Q(\core.CPU_Dmem_value_a5[10][31] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][3]$_SDFFE_PP1P_  (.D(_00265_),
    .Q(\core.CPU_Dmem_value_a5[10][3] ),
    .CLK(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][4]$_SDFFE_PP0P_  (.D(_00266_),
    .Q(\core.CPU_Dmem_value_a5[10][4] ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][5]$_SDFFE_PP0P_  (.D(_00267_),
    .Q(\core.CPU_Dmem_value_a5[10][5] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][6]$_SDFFE_PP0P_  (.D(_00268_),
    .Q(\core.CPU_Dmem_value_a5[10][6] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][7]$_SDFFE_PP0P_  (.D(_00269_),
    .Q(\core.CPU_Dmem_value_a5[10][7] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][8]$_SDFFE_PP0P_  (.D(_00270_),
    .Q(\core.CPU_Dmem_value_a5[10][8] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[10][9]$_SDFFE_PP0P_  (.D(_00271_),
    .Q(\core.CPU_Dmem_value_a5[10][9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][0]$_SDFFE_PP1P_  (.D(_00272_),
    .Q(\core.CPU_Dmem_value_a5[11][0] ),
    .CLK(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][10]$_SDFFE_PP0P_  (.D(_00273_),
    .Q(\core.CPU_Dmem_value_a5[11][10] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][11]$_SDFFE_PP0P_  (.D(_00274_),
    .Q(\core.CPU_Dmem_value_a5[11][11] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][12]$_SDFFE_PP0P_  (.D(_00275_),
    .Q(\core.CPU_Dmem_value_a5[11][12] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][13]$_SDFFE_PP0P_  (.D(_00276_),
    .Q(\core.CPU_Dmem_value_a5[11][13] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][14]$_SDFFE_PP0P_  (.D(_00277_),
    .Q(\core.CPU_Dmem_value_a5[11][14] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][15]$_SDFFE_PP0P_  (.D(_00278_),
    .Q(\core.CPU_Dmem_value_a5[11][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][16]$_SDFFE_PP0P_  (.D(_00279_),
    .Q(\core.CPU_Dmem_value_a5[11][16] ),
    .CLK(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][17]$_SDFFE_PP0P_  (.D(_00280_),
    .Q(\core.CPU_Dmem_value_a5[11][17] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][18]$_SDFFE_PP0P_  (.D(_00281_),
    .Q(\core.CPU_Dmem_value_a5[11][18] ),
    .CLK(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][19]$_SDFFE_PP0P_  (.D(_00282_),
    .Q(\core.CPU_Dmem_value_a5[11][19] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][1]$_SDFFE_PP1P_  (.D(_00283_),
    .Q(\core.CPU_Dmem_value_a5[11][1] ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][20]$_SDFFE_PP0P_  (.D(_00284_),
    .Q(\core.CPU_Dmem_value_a5[11][20] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][21]$_SDFFE_PP0P_  (.D(_00285_),
    .Q(\core.CPU_Dmem_value_a5[11][21] ),
    .CLK(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][22]$_SDFFE_PP0P_  (.D(_00286_),
    .Q(\core.CPU_Dmem_value_a5[11][22] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][23]$_SDFFE_PP0P_  (.D(_00287_),
    .Q(\core.CPU_Dmem_value_a5[11][23] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][24]$_SDFFE_PP0P_  (.D(_00288_),
    .Q(\core.CPU_Dmem_value_a5[11][24] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][25]$_SDFFE_PP0P_  (.D(_00289_),
    .Q(\core.CPU_Dmem_value_a5[11][25] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][26]$_SDFFE_PP0P_  (.D(_00290_),
    .Q(\core.CPU_Dmem_value_a5[11][26] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][27]$_SDFFE_PP0P_  (.D(_00291_),
    .Q(\core.CPU_Dmem_value_a5[11][27] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][28]$_SDFFE_PP0P_  (.D(_00292_),
    .Q(\core.CPU_Dmem_value_a5[11][28] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][29]$_SDFFE_PP0P_  (.D(_00293_),
    .Q(\core.CPU_Dmem_value_a5[11][29] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][2]$_SDFFE_PP0P_  (.D(_00294_),
    .Q(\core.CPU_Dmem_value_a5[11][2] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][30]$_SDFFE_PP0P_  (.D(_00295_),
    .Q(\core.CPU_Dmem_value_a5[11][30] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][31]$_SDFFE_PP0P_  (.D(_00296_),
    .Q(\core.CPU_Dmem_value_a5[11][31] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][3]$_SDFFE_PP1P_  (.D(_00297_),
    .Q(\core.CPU_Dmem_value_a5[11][3] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][4]$_SDFFE_PP0P_  (.D(_00298_),
    .Q(\core.CPU_Dmem_value_a5[11][4] ),
    .CLK(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][5]$_SDFFE_PP0P_  (.D(_00299_),
    .Q(\core.CPU_Dmem_value_a5[11][5] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][6]$_SDFFE_PP0P_  (.D(_00300_),
    .Q(\core.CPU_Dmem_value_a5[11][6] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][7]$_SDFFE_PP0P_  (.D(_00301_),
    .Q(\core.CPU_Dmem_value_a5[11][7] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][8]$_SDFFE_PP0P_  (.D(_00302_),
    .Q(\core.CPU_Dmem_value_a5[11][8] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[11][9]$_SDFFE_PP0P_  (.D(_00303_),
    .Q(\core.CPU_Dmem_value_a5[11][9] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][0]$_SDFFE_PP0P_  (.D(_00304_),
    .Q(\core.CPU_Dmem_value_a5[12][0] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][10]$_SDFFE_PP0P_  (.D(_00305_),
    .Q(\core.CPU_Dmem_value_a5[12][10] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][11]$_SDFFE_PP0P_  (.D(_00306_),
    .Q(\core.CPU_Dmem_value_a5[12][11] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][12]$_SDFFE_PP0P_  (.D(_00307_),
    .Q(\core.CPU_Dmem_value_a5[12][12] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][13]$_SDFFE_PP0P_  (.D(_00308_),
    .Q(\core.CPU_Dmem_value_a5[12][13] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][14]$_SDFFE_PP0P_  (.D(_00309_),
    .Q(\core.CPU_Dmem_value_a5[12][14] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][15]$_SDFFE_PP0P_  (.D(_00310_),
    .Q(\core.CPU_Dmem_value_a5[12][15] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][16]$_SDFFE_PP0P_  (.D(_00311_),
    .Q(\core.CPU_Dmem_value_a5[12][16] ),
    .CLK(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][17]$_SDFFE_PP0P_  (.D(_00312_),
    .Q(\core.CPU_Dmem_value_a5[12][17] ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][18]$_SDFFE_PP0P_  (.D(_00313_),
    .Q(\core.CPU_Dmem_value_a5[12][18] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][19]$_SDFFE_PP0P_  (.D(_00314_),
    .Q(\core.CPU_Dmem_value_a5[12][19] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][1]$_SDFFE_PP0P_  (.D(_00315_),
    .Q(\core.CPU_Dmem_value_a5[12][1] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][20]$_SDFFE_PP0P_  (.D(_00316_),
    .Q(\core.CPU_Dmem_value_a5[12][20] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][21]$_SDFFE_PP0P_  (.D(_00317_),
    .Q(\core.CPU_Dmem_value_a5[12][21] ),
    .CLK(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][22]$_SDFFE_PP0P_  (.D(_00318_),
    .Q(\core.CPU_Dmem_value_a5[12][22] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][23]$_SDFFE_PP0P_  (.D(_00319_),
    .Q(\core.CPU_Dmem_value_a5[12][23] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][24]$_SDFFE_PP0P_  (.D(_00320_),
    .Q(\core.CPU_Dmem_value_a5[12][24] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][25]$_SDFFE_PP0P_  (.D(_00321_),
    .Q(\core.CPU_Dmem_value_a5[12][25] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][26]$_SDFFE_PP0P_  (.D(_00322_),
    .Q(\core.CPU_Dmem_value_a5[12][26] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][27]$_SDFFE_PP0P_  (.D(_00323_),
    .Q(\core.CPU_Dmem_value_a5[12][27] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][28]$_SDFFE_PP0P_  (.D(_00324_),
    .Q(\core.CPU_Dmem_value_a5[12][28] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][29]$_SDFFE_PP0P_  (.D(_00325_),
    .Q(\core.CPU_Dmem_value_a5[12][29] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][2]$_SDFFE_PP1P_  (.D(_00326_),
    .Q(\core.CPU_Dmem_value_a5[12][2] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][30]$_SDFFE_PP0P_  (.D(_00327_),
    .Q(\core.CPU_Dmem_value_a5[12][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][31]$_SDFFE_PP0P_  (.D(_00328_),
    .Q(\core.CPU_Dmem_value_a5[12][31] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][3]$_SDFFE_PP1P_  (.D(_00329_),
    .Q(\core.CPU_Dmem_value_a5[12][3] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][4]$_SDFFE_PP0P_  (.D(_00330_),
    .Q(\core.CPU_Dmem_value_a5[12][4] ),
    .CLK(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][5]$_SDFFE_PP0P_  (.D(_00331_),
    .Q(\core.CPU_Dmem_value_a5[12][5] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][6]$_SDFFE_PP0P_  (.D(_00332_),
    .Q(\core.CPU_Dmem_value_a5[12][6] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][7]$_SDFFE_PP0P_  (.D(_00333_),
    .Q(\core.CPU_Dmem_value_a5[12][7] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][8]$_SDFFE_PP0P_  (.D(_00334_),
    .Q(\core.CPU_Dmem_value_a5[12][8] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[12][9]$_SDFFE_PP0P_  (.D(_00335_),
    .Q(\core.CPU_Dmem_value_a5[12][9] ),
    .CLK(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][0]$_SDFFE_PP1P_  (.D(_00336_),
    .Q(\core.CPU_Dmem_value_a5[13][0] ),
    .CLK(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][10]$_SDFFE_PP0P_  (.D(_00337_),
    .Q(\core.CPU_Dmem_value_a5[13][10] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][11]$_SDFFE_PP0P_  (.D(_00338_),
    .Q(\core.CPU_Dmem_value_a5[13][11] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][12]$_SDFFE_PP0P_  (.D(_00339_),
    .Q(\core.CPU_Dmem_value_a5[13][12] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][13]$_SDFFE_PP0P_  (.D(_00340_),
    .Q(\core.CPU_Dmem_value_a5[13][13] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][14]$_SDFFE_PP0P_  (.D(_00341_),
    .Q(\core.CPU_Dmem_value_a5[13][14] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][15]$_SDFFE_PP0P_  (.D(_00342_),
    .Q(\core.CPU_Dmem_value_a5[13][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][16]$_SDFFE_PP0P_  (.D(_00343_),
    .Q(\core.CPU_Dmem_value_a5[13][16] ),
    .CLK(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][17]$_SDFFE_PP0P_  (.D(_00344_),
    .Q(\core.CPU_Dmem_value_a5[13][17] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][18]$_SDFFE_PP0P_  (.D(_00345_),
    .Q(\core.CPU_Dmem_value_a5[13][18] ),
    .CLK(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][19]$_SDFFE_PP0P_  (.D(_00346_),
    .Q(\core.CPU_Dmem_value_a5[13][19] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][1]$_SDFFE_PP0P_  (.D(_00347_),
    .Q(\core.CPU_Dmem_value_a5[13][1] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][20]$_SDFFE_PP0P_  (.D(_00348_),
    .Q(\core.CPU_Dmem_value_a5[13][20] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][21]$_SDFFE_PP0P_  (.D(_00349_),
    .Q(\core.CPU_Dmem_value_a5[13][21] ),
    .CLK(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][22]$_SDFFE_PP0P_  (.D(_00350_),
    .Q(\core.CPU_Dmem_value_a5[13][22] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][23]$_SDFFE_PP0P_  (.D(_00351_),
    .Q(\core.CPU_Dmem_value_a5[13][23] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][24]$_SDFFE_PP0P_  (.D(_00352_),
    .Q(\core.CPU_Dmem_value_a5[13][24] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][25]$_SDFFE_PP0P_  (.D(_00353_),
    .Q(\core.CPU_Dmem_value_a5[13][25] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][26]$_SDFFE_PP0P_  (.D(_00354_),
    .Q(\core.CPU_Dmem_value_a5[13][26] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][27]$_SDFFE_PP0P_  (.D(_00355_),
    .Q(\core.CPU_Dmem_value_a5[13][27] ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][28]$_SDFFE_PP0P_  (.D(_00356_),
    .Q(\core.CPU_Dmem_value_a5[13][28] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][29]$_SDFFE_PP0P_  (.D(_00357_),
    .Q(\core.CPU_Dmem_value_a5[13][29] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][2]$_SDFFE_PP1P_  (.D(_00358_),
    .Q(\core.CPU_Dmem_value_a5[13][2] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][30]$_SDFFE_PP0P_  (.D(_00359_),
    .Q(\core.CPU_Dmem_value_a5[13][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][31]$_SDFFE_PP0P_  (.D(_00360_),
    .Q(\core.CPU_Dmem_value_a5[13][31] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][3]$_SDFFE_PP1P_  (.D(_00361_),
    .Q(\core.CPU_Dmem_value_a5[13][3] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][4]$_SDFFE_PP0P_  (.D(_00362_),
    .Q(\core.CPU_Dmem_value_a5[13][4] ),
    .CLK(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][5]$_SDFFE_PP0P_  (.D(_00363_),
    .Q(\core.CPU_Dmem_value_a5[13][5] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][6]$_SDFFE_PP0P_  (.D(_00364_),
    .Q(\core.CPU_Dmem_value_a5[13][6] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][7]$_SDFFE_PP0P_  (.D(_00365_),
    .Q(\core.CPU_Dmem_value_a5[13][7] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][8]$_SDFFE_PP0P_  (.D(_00366_),
    .Q(\core.CPU_Dmem_value_a5[13][8] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[13][9]$_SDFFE_PP0P_  (.D(_00367_),
    .Q(\core.CPU_Dmem_value_a5[13][9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][0]$_SDFFE_PP0P_  (.D(_00368_),
    .Q(\core.CPU_Dmem_value_a5[14][0] ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][10]$_SDFFE_PP0P_  (.D(_00369_),
    .Q(\core.CPU_Dmem_value_a5[14][10] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][11]$_SDFFE_PP0P_  (.D(_00370_),
    .Q(\core.CPU_Dmem_value_a5[14][11] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][12]$_SDFFE_PP0P_  (.D(_00371_),
    .Q(\core.CPU_Dmem_value_a5[14][12] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][13]$_SDFFE_PP0P_  (.D(_00372_),
    .Q(\core.CPU_Dmem_value_a5[14][13] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][14]$_SDFFE_PP0P_  (.D(_00373_),
    .Q(\core.CPU_Dmem_value_a5[14][14] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][15]$_SDFFE_PP0P_  (.D(_00374_),
    .Q(\core.CPU_Dmem_value_a5[14][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][16]$_SDFFE_PP0P_  (.D(_00375_),
    .Q(\core.CPU_Dmem_value_a5[14][16] ),
    .CLK(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][17]$_SDFFE_PP0P_  (.D(_00376_),
    .Q(\core.CPU_Dmem_value_a5[14][17] ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][18]$_SDFFE_PP0P_  (.D(_00377_),
    .Q(\core.CPU_Dmem_value_a5[14][18] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][19]$_SDFFE_PP0P_  (.D(_00378_),
    .Q(\core.CPU_Dmem_value_a5[14][19] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][1]$_SDFFE_PP1P_  (.D(_00379_),
    .Q(\core.CPU_Dmem_value_a5[14][1] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][20]$_SDFFE_PP0P_  (.D(_00380_),
    .Q(\core.CPU_Dmem_value_a5[14][20] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][21]$_SDFFE_PP0P_  (.D(_00381_),
    .Q(\core.CPU_Dmem_value_a5[14][21] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][22]$_SDFFE_PP0P_  (.D(_00382_),
    .Q(\core.CPU_Dmem_value_a5[14][22] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][23]$_SDFFE_PP0P_  (.D(_00383_),
    .Q(\core.CPU_Dmem_value_a5[14][23] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][24]$_SDFFE_PP0P_  (.D(_00384_),
    .Q(\core.CPU_Dmem_value_a5[14][24] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][25]$_SDFFE_PP0P_  (.D(_00385_),
    .Q(\core.CPU_Dmem_value_a5[14][25] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][26]$_SDFFE_PP0P_  (.D(_00386_),
    .Q(\core.CPU_Dmem_value_a5[14][26] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][27]$_SDFFE_PP0P_  (.D(_00387_),
    .Q(\core.CPU_Dmem_value_a5[14][27] ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][28]$_SDFFE_PP0P_  (.D(_00388_),
    .Q(\core.CPU_Dmem_value_a5[14][28] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][29]$_SDFFE_PP0P_  (.D(_00389_),
    .Q(\core.CPU_Dmem_value_a5[14][29] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][2]$_SDFFE_PP1P_  (.D(_00390_),
    .Q(\core.CPU_Dmem_value_a5[14][2] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][30]$_SDFFE_PP0P_  (.D(_00391_),
    .Q(\core.CPU_Dmem_value_a5[14][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][31]$_SDFFE_PP0P_  (.D(_00392_),
    .Q(\core.CPU_Dmem_value_a5[14][31] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][3]$_SDFFE_PP1P_  (.D(_00393_),
    .Q(\core.CPU_Dmem_value_a5[14][3] ),
    .CLK(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][4]$_SDFFE_PP0P_  (.D(_00394_),
    .Q(\core.CPU_Dmem_value_a5[14][4] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][5]$_SDFFE_PP0P_  (.D(_00395_),
    .Q(\core.CPU_Dmem_value_a5[14][5] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][6]$_SDFFE_PP0P_  (.D(_00396_),
    .Q(\core.CPU_Dmem_value_a5[14][6] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][7]$_SDFFE_PP0P_  (.D(_00397_),
    .Q(\core.CPU_Dmem_value_a5[14][7] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][8]$_SDFFE_PP0P_  (.D(_00398_),
    .Q(\core.CPU_Dmem_value_a5[14][8] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[14][9]$_SDFFE_PP0P_  (.D(_00399_),
    .Q(\core.CPU_Dmem_value_a5[14][9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][0]$_SDFFE_PP1P_  (.D(_00400_),
    .Q(\core.CPU_Dmem_value_a5[15][0] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][10]$_SDFFE_PP0P_  (.D(_00401_),
    .Q(\core.CPU_Dmem_value_a5[15][10] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][11]$_SDFFE_PP0P_  (.D(_00402_),
    .Q(\core.CPU_Dmem_value_a5[15][11] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][12]$_SDFFE_PP0P_  (.D(_00403_),
    .Q(\core.CPU_Dmem_value_a5[15][12] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][13]$_SDFFE_PP0P_  (.D(_00404_),
    .Q(\core.CPU_Dmem_value_a5[15][13] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][14]$_SDFFE_PP0P_  (.D(_00405_),
    .Q(\core.CPU_Dmem_value_a5[15][14] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][15]$_SDFFE_PP0P_  (.D(_00406_),
    .Q(\core.CPU_Dmem_value_a5[15][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][16]$_SDFFE_PP0P_  (.D(_00407_),
    .Q(\core.CPU_Dmem_value_a5[15][16] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][17]$_SDFFE_PP0P_  (.D(_00408_),
    .Q(\core.CPU_Dmem_value_a5[15][17] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][18]$_SDFFE_PP0P_  (.D(_00409_),
    .Q(\core.CPU_Dmem_value_a5[15][18] ),
    .CLK(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][19]$_SDFFE_PP0P_  (.D(_00410_),
    .Q(\core.CPU_Dmem_value_a5[15][19] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][1]$_SDFFE_PP1P_  (.D(_00411_),
    .Q(\core.CPU_Dmem_value_a5[15][1] ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][20]$_SDFFE_PP0P_  (.D(_00412_),
    .Q(\core.CPU_Dmem_value_a5[15][20] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][21]$_SDFFE_PP0P_  (.D(_00413_),
    .Q(\core.CPU_Dmem_value_a5[15][21] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][22]$_SDFFE_PP0P_  (.D(_00414_),
    .Q(\core.CPU_Dmem_value_a5[15][22] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][23]$_SDFFE_PP0P_  (.D(_00415_),
    .Q(\core.CPU_Dmem_value_a5[15][23] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][24]$_SDFFE_PP0P_  (.D(_00416_),
    .Q(\core.CPU_Dmem_value_a5[15][24] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][25]$_SDFFE_PP0P_  (.D(_00417_),
    .Q(\core.CPU_Dmem_value_a5[15][25] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][26]$_SDFFE_PP0P_  (.D(_00418_),
    .Q(\core.CPU_Dmem_value_a5[15][26] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][27]$_SDFFE_PP0P_  (.D(_00419_),
    .Q(\core.CPU_Dmem_value_a5[15][27] ),
    .CLK(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][28]$_SDFFE_PP0P_  (.D(_00420_),
    .Q(\core.CPU_Dmem_value_a5[15][28] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][29]$_SDFFE_PP0P_  (.D(_00421_),
    .Q(\core.CPU_Dmem_value_a5[15][29] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][2]$_SDFFE_PP1P_  (.D(_00422_),
    .Q(\core.CPU_Dmem_value_a5[15][2] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][30]$_SDFFE_PP0P_  (.D(_00423_),
    .Q(\core.CPU_Dmem_value_a5[15][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][31]$_SDFFE_PP0P_  (.D(_00424_),
    .Q(\core.CPU_Dmem_value_a5[15][31] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][3]$_SDFFE_PP1P_  (.D(_00425_),
    .Q(\core.CPU_Dmem_value_a5[15][3] ),
    .CLK(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][4]$_SDFFE_PP0P_  (.D(_00426_),
    .Q(\core.CPU_Dmem_value_a5[15][4] ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][5]$_SDFFE_PP0P_  (.D(_00427_),
    .Q(\core.CPU_Dmem_value_a5[15][5] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][6]$_SDFFE_PP0P_  (.D(_00428_),
    .Q(\core.CPU_Dmem_value_a5[15][6] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][7]$_SDFFE_PP0P_  (.D(_00429_),
    .Q(\core.CPU_Dmem_value_a5[15][7] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][8]$_SDFFE_PP0P_  (.D(_00430_),
    .Q(\core.CPU_Dmem_value_a5[15][8] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[15][9]$_SDFFE_PP0P_  (.D(_00431_),
    .Q(\core.CPU_Dmem_value_a5[15][9] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][0]$_SDFFE_PP1P_  (.D(_00432_),
    .Q(\core.CPU_Dmem_value_a5[1][0] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][10]$_SDFFE_PP0P_  (.D(_00433_),
    .Q(\core.CPU_Dmem_value_a5[1][10] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][11]$_SDFFE_PP0P_  (.D(_00434_),
    .Q(\core.CPU_Dmem_value_a5[1][11] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][12]$_SDFFE_PP0P_  (.D(_00435_),
    .Q(\core.CPU_Dmem_value_a5[1][12] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][13]$_SDFFE_PP0P_  (.D(_00436_),
    .Q(\core.CPU_Dmem_value_a5[1][13] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][14]$_SDFFE_PP0P_  (.D(_00437_),
    .Q(\core.CPU_Dmem_value_a5[1][14] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][15]$_SDFFE_PP0P_  (.D(_00438_),
    .Q(\core.CPU_Dmem_value_a5[1][15] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][16]$_SDFFE_PP0P_  (.D(_00439_),
    .Q(\core.CPU_Dmem_value_a5[1][16] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][17]$_SDFFE_PP0P_  (.D(_00440_),
    .Q(\core.CPU_Dmem_value_a5[1][17] ),
    .CLK(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][18]$_SDFFE_PP0P_  (.D(_00441_),
    .Q(\core.CPU_Dmem_value_a5[1][18] ),
    .CLK(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][19]$_SDFFE_PP0P_  (.D(_00442_),
    .Q(\core.CPU_Dmem_value_a5[1][19] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][1]$_SDFFE_PP0P_  (.D(_00443_),
    .Q(\core.CPU_Dmem_value_a5[1][1] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][20]$_SDFFE_PP0P_  (.D(_00444_),
    .Q(\core.CPU_Dmem_value_a5[1][20] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][21]$_SDFFE_PP0P_  (.D(_00445_),
    .Q(\core.CPU_Dmem_value_a5[1][21] ),
    .CLK(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][22]$_SDFFE_PP0P_  (.D(_00446_),
    .Q(\core.CPU_Dmem_value_a5[1][22] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][23]$_SDFFE_PP0P_  (.D(_00447_),
    .Q(\core.CPU_Dmem_value_a5[1][23] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][24]$_SDFFE_PP0P_  (.D(_00448_),
    .Q(\core.CPU_Dmem_value_a5[1][24] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][25]$_SDFFE_PP0P_  (.D(_00449_),
    .Q(\core.CPU_Dmem_value_a5[1][25] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][26]$_SDFFE_PP0P_  (.D(_00450_),
    .Q(\core.CPU_Dmem_value_a5[1][26] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][27]$_SDFFE_PP0P_  (.D(_00451_),
    .Q(\core.CPU_Dmem_value_a5[1][27] ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][28]$_SDFFE_PP0P_  (.D(_00452_),
    .Q(\core.CPU_Dmem_value_a5[1][28] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][29]$_SDFFE_PP0P_  (.D(_00453_),
    .Q(\core.CPU_Dmem_value_a5[1][29] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][2]$_SDFFE_PP0P_  (.D(_00454_),
    .Q(\core.CPU_Dmem_value_a5[1][2] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][30]$_SDFFE_PP0P_  (.D(_00455_),
    .Q(\core.CPU_Dmem_value_a5[1][30] ),
    .CLK(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][31]$_SDFFE_PP0P_  (.D(_00456_),
    .Q(\core.CPU_Dmem_value_a5[1][31] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][3]$_SDFFE_PP0P_  (.D(_00457_),
    .Q(\core.CPU_Dmem_value_a5[1][3] ),
    .CLK(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][4]$_SDFFE_PP0P_  (.D(_00458_),
    .Q(\core.CPU_Dmem_value_a5[1][4] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][5]$_SDFFE_PP0P_  (.D(_00459_),
    .Q(\core.CPU_Dmem_value_a5[1][5] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][6]$_SDFFE_PP0P_  (.D(_00460_),
    .Q(\core.CPU_Dmem_value_a5[1][6] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][7]$_SDFFE_PP0P_  (.D(_00461_),
    .Q(\core.CPU_Dmem_value_a5[1][7] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][8]$_SDFFE_PP0P_  (.D(_00462_),
    .Q(\core.CPU_Dmem_value_a5[1][8] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[1][9]$_SDFFE_PP0P_  (.D(_00463_),
    .Q(\core.CPU_Dmem_value_a5[1][9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][0]$_SDFFE_PP0P_  (.D(_00464_),
    .Q(\core.CPU_Dmem_value_a5[2][0] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][10]$_SDFFE_PP0P_  (.D(_00465_),
    .Q(\core.CPU_Dmem_value_a5[2][10] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][11]$_SDFFE_PP0P_  (.D(_00466_),
    .Q(\core.CPU_Dmem_value_a5[2][11] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][12]$_SDFFE_PP0P_  (.D(_00467_),
    .Q(\core.CPU_Dmem_value_a5[2][12] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][13]$_SDFFE_PP0P_  (.D(_00468_),
    .Q(\core.CPU_Dmem_value_a5[2][13] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][14]$_SDFFE_PP0P_  (.D(_00469_),
    .Q(\core.CPU_Dmem_value_a5[2][14] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][15]$_SDFFE_PP0P_  (.D(_00470_),
    .Q(\core.CPU_Dmem_value_a5[2][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][16]$_SDFFE_PP0P_  (.D(_00471_),
    .Q(\core.CPU_Dmem_value_a5[2][16] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][17]$_SDFFE_PP0P_  (.D(_00472_),
    .Q(\core.CPU_Dmem_value_a5[2][17] ),
    .CLK(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][18]$_SDFFE_PP0P_  (.D(_00473_),
    .Q(\core.CPU_Dmem_value_a5[2][18] ),
    .CLK(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][19]$_SDFFE_PP0P_  (.D(_00474_),
    .Q(\core.CPU_Dmem_value_a5[2][19] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][1]$_SDFFE_PP1P_  (.D(_00475_),
    .Q(\core.CPU_Dmem_value_a5[2][1] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][20]$_SDFFE_PP0P_  (.D(_00476_),
    .Q(\core.CPU_Dmem_value_a5[2][20] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][21]$_SDFFE_PP0P_  (.D(_00477_),
    .Q(\core.CPU_Dmem_value_a5[2][21] ),
    .CLK(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][22]$_SDFFE_PP0P_  (.D(_00478_),
    .Q(\core.CPU_Dmem_value_a5[2][22] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][23]$_SDFFE_PP0P_  (.D(_00479_),
    .Q(\core.CPU_Dmem_value_a5[2][23] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][24]$_SDFFE_PP0P_  (.D(_00480_),
    .Q(\core.CPU_Dmem_value_a5[2][24] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][25]$_SDFFE_PP0P_  (.D(_00481_),
    .Q(\core.CPU_Dmem_value_a5[2][25] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][26]$_SDFFE_PP0P_  (.D(_00482_),
    .Q(\core.CPU_Dmem_value_a5[2][26] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][27]$_SDFFE_PP0P_  (.D(_00483_),
    .Q(\core.CPU_Dmem_value_a5[2][27] ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][28]$_SDFFE_PP0P_  (.D(_00484_),
    .Q(\core.CPU_Dmem_value_a5[2][28] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][29]$_SDFFE_PP0P_  (.D(_00485_),
    .Q(\core.CPU_Dmem_value_a5[2][29] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][2]$_SDFFE_PP0P_  (.D(_00486_),
    .Q(\core.CPU_Dmem_value_a5[2][2] ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][30]$_SDFFE_PP0P_  (.D(_00487_),
    .Q(\core.CPU_Dmem_value_a5[2][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][31]$_SDFFE_PP0P_  (.D(_00488_),
    .Q(\core.CPU_Dmem_value_a5[2][31] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][3]$_SDFFE_PP0P_  (.D(_00489_),
    .Q(\core.CPU_Dmem_value_a5[2][3] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][4]$_SDFFE_PP0P_  (.D(_00490_),
    .Q(\core.CPU_Dmem_value_a5[2][4] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][5]$_SDFFE_PP0P_  (.D(_00491_),
    .Q(\core.CPU_Dmem_value_a5[2][5] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][6]$_SDFFE_PP0P_  (.D(_00492_),
    .Q(\core.CPU_Dmem_value_a5[2][6] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][7]$_SDFFE_PP0P_  (.D(_00493_),
    .Q(\core.CPU_Dmem_value_a5[2][7] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][8]$_SDFFE_PP0P_  (.D(_00494_),
    .Q(\core.CPU_Dmem_value_a5[2][8] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[2][9]$_SDFFE_PP0P_  (.D(_00495_),
    .Q(\core.CPU_Dmem_value_a5[2][9] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][0]$_SDFFE_PP1P_  (.D(_00496_),
    .Q(\core.CPU_Dmem_value_a5[3][0] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][10]$_SDFFE_PP0P_  (.D(_00497_),
    .Q(\core.CPU_Dmem_value_a5[3][10] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][11]$_SDFFE_PP0P_  (.D(_00498_),
    .Q(\core.CPU_Dmem_value_a5[3][11] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][12]$_SDFFE_PP0P_  (.D(_00499_),
    .Q(\core.CPU_Dmem_value_a5[3][12] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][13]$_SDFFE_PP0P_  (.D(_00500_),
    .Q(\core.CPU_Dmem_value_a5[3][13] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][14]$_SDFFE_PP0P_  (.D(_00501_),
    .Q(\core.CPU_Dmem_value_a5[3][14] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][15]$_SDFFE_PP0P_  (.D(_00502_),
    .Q(\core.CPU_Dmem_value_a5[3][15] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][16]$_SDFFE_PP0P_  (.D(_00503_),
    .Q(\core.CPU_Dmem_value_a5[3][16] ),
    .CLK(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][17]$_SDFFE_PP0P_  (.D(_00504_),
    .Q(\core.CPU_Dmem_value_a5[3][17] ),
    .CLK(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][18]$_SDFFE_PP0P_  (.D(_00505_),
    .Q(\core.CPU_Dmem_value_a5[3][18] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][19]$_SDFFE_PP0P_  (.D(_00506_),
    .Q(\core.CPU_Dmem_value_a5[3][19] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][1]$_SDFFE_PP1P_  (.D(_00507_),
    .Q(\core.CPU_Dmem_value_a5[3][1] ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][20]$_SDFFE_PP0P_  (.D(_00508_),
    .Q(\core.CPU_Dmem_value_a5[3][20] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][21]$_SDFFE_PP0P_  (.D(_00509_),
    .Q(\core.CPU_Dmem_value_a5[3][21] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][22]$_SDFFE_PP0P_  (.D(_00510_),
    .Q(\core.CPU_Dmem_value_a5[3][22] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][23]$_SDFFE_PP0P_  (.D(_00511_),
    .Q(\core.CPU_Dmem_value_a5[3][23] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][24]$_SDFFE_PP0P_  (.D(_00512_),
    .Q(\core.CPU_Dmem_value_a5[3][24] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][25]$_SDFFE_PP0P_  (.D(_00513_),
    .Q(\core.CPU_Dmem_value_a5[3][25] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][26]$_SDFFE_PP0P_  (.D(_00514_),
    .Q(\core.CPU_Dmem_value_a5[3][26] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][27]$_SDFFE_PP0P_  (.D(_00515_),
    .Q(\core.CPU_Dmem_value_a5[3][27] ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][28]$_SDFFE_PP0P_  (.D(_00516_),
    .Q(\core.CPU_Dmem_value_a5[3][28] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][29]$_SDFFE_PP0P_  (.D(_00517_),
    .Q(\core.CPU_Dmem_value_a5[3][29] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][2]$_SDFFE_PP0P_  (.D(_00518_),
    .Q(\core.CPU_Dmem_value_a5[3][2] ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][30]$_SDFFE_PP0P_  (.D(_00519_),
    .Q(\core.CPU_Dmem_value_a5[3][30] ),
    .CLK(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][31]$_SDFFE_PP0P_  (.D(_00520_),
    .Q(\core.CPU_Dmem_value_a5[3][31] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][3]$_SDFFE_PP0P_  (.D(_00521_),
    .Q(\core.CPU_Dmem_value_a5[3][3] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][4]$_SDFFE_PP0P_  (.D(_00522_),
    .Q(\core.CPU_Dmem_value_a5[3][4] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][5]$_SDFFE_PP0P_  (.D(_00523_),
    .Q(\core.CPU_Dmem_value_a5[3][5] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][6]$_SDFFE_PP0P_  (.D(_00524_),
    .Q(\core.CPU_Dmem_value_a5[3][6] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][7]$_SDFFE_PP0P_  (.D(_00525_),
    .Q(\core.CPU_Dmem_value_a5[3][7] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][8]$_SDFFE_PP0P_  (.D(_00526_),
    .Q(\core.CPU_Dmem_value_a5[3][8] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[3][9]$_SDFFE_PP0P_  (.D(_00527_),
    .Q(\core.CPU_Dmem_value_a5[3][9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][0]$_SDFFE_PP0P_  (.D(_00528_),
    .Q(\core.CPU_Dmem_value_a5[4][0] ),
    .CLK(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][10]$_SDFFE_PP0P_  (.D(_00529_),
    .Q(\core.CPU_Dmem_value_a5[4][10] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][11]$_SDFFE_PP0P_  (.D(_00530_),
    .Q(\core.CPU_Dmem_value_a5[4][11] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][12]$_SDFFE_PP0P_  (.D(_00531_),
    .Q(\core.CPU_Dmem_value_a5[4][12] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][13]$_SDFFE_PP0P_  (.D(_00532_),
    .Q(\core.CPU_Dmem_value_a5[4][13] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][14]$_SDFFE_PP0P_  (.D(_00533_),
    .Q(\core.CPU_Dmem_value_a5[4][14] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][15]$_SDFFE_PP0P_  (.D(_00534_),
    .Q(\core.CPU_Dmem_value_a5[4][15] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][16]$_SDFFE_PP0P_  (.D(_00535_),
    .Q(\core.CPU_Dmem_value_a5[4][16] ),
    .CLK(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][17]$_SDFFE_PP0P_  (.D(_00536_),
    .Q(\core.CPU_Dmem_value_a5[4][17] ),
    .CLK(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][18]$_SDFFE_PP0P_  (.D(_00537_),
    .Q(\core.CPU_Dmem_value_a5[4][18] ),
    .CLK(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][19]$_SDFFE_PP0P_  (.D(_00538_),
    .Q(\core.CPU_Dmem_value_a5[4][19] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][1]$_SDFFE_PP0P_  (.D(_00539_),
    .Q(\core.CPU_Dmem_value_a5[4][1] ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][20]$_SDFFE_PP0P_  (.D(_00540_),
    .Q(\core.CPU_Dmem_value_a5[4][20] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][21]$_SDFFE_PP0P_  (.D(_00541_),
    .Q(\core.CPU_Dmem_value_a5[4][21] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][22]$_SDFFE_PP0P_  (.D(_00542_),
    .Q(\core.CPU_Dmem_value_a5[4][22] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][23]$_SDFFE_PP0P_  (.D(_00543_),
    .Q(\core.CPU_Dmem_value_a5[4][23] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][24]$_SDFFE_PP0P_  (.D(_00544_),
    .Q(\core.CPU_Dmem_value_a5[4][24] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][25]$_SDFFE_PP0P_  (.D(_00545_),
    .Q(\core.CPU_Dmem_value_a5[4][25] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][26]$_SDFFE_PP0P_  (.D(_00546_),
    .Q(\core.CPU_Dmem_value_a5[4][26] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][27]$_SDFFE_PP0P_  (.D(_00547_),
    .Q(\core.CPU_Dmem_value_a5[4][27] ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][28]$_SDFFE_PP0P_  (.D(_00548_),
    .Q(\core.CPU_Dmem_value_a5[4][28] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][29]$_SDFFE_PP0P_  (.D(_00549_),
    .Q(\core.CPU_Dmem_value_a5[4][29] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][2]$_SDFFE_PP1P_  (.D(_00550_),
    .Q(\core.CPU_Dmem_value_a5[4][2] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][30]$_SDFFE_PP0P_  (.D(_00551_),
    .Q(\core.CPU_Dmem_value_a5[4][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][31]$_SDFFE_PP0P_  (.D(_00552_),
    .Q(\core.CPU_Dmem_value_a5[4][31] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][3]$_SDFFE_PP0P_  (.D(_00553_),
    .Q(\core.CPU_Dmem_value_a5[4][3] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][4]$_SDFFE_PP0P_  (.D(_00554_),
    .Q(\core.CPU_Dmem_value_a5[4][4] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][5]$_SDFFE_PP0P_  (.D(_00555_),
    .Q(\core.CPU_Dmem_value_a5[4][5] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][6]$_SDFFE_PP0P_  (.D(_00556_),
    .Q(\core.CPU_Dmem_value_a5[4][6] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][7]$_SDFFE_PP0P_  (.D(_00557_),
    .Q(\core.CPU_Dmem_value_a5[4][7] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][8]$_SDFFE_PP0P_  (.D(_00558_),
    .Q(\core.CPU_Dmem_value_a5[4][8] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[4][9]$_SDFFE_PP0P_  (.D(_00559_),
    .Q(\core.CPU_Dmem_value_a5[4][9] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][0]$_SDFFE_PP1P_  (.D(_00560_),
    .Q(\core.CPU_Dmem_value_a5[5][0] ),
    .CLK(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][10]$_SDFFE_PP0P_  (.D(_00561_),
    .Q(\core.CPU_Dmem_value_a5[5][10] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][11]$_SDFFE_PP0P_  (.D(_00562_),
    .Q(\core.CPU_Dmem_value_a5[5][11] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][12]$_SDFFE_PP0P_  (.D(_00563_),
    .Q(\core.CPU_Dmem_value_a5[5][12] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][13]$_SDFFE_PP0P_  (.D(_00564_),
    .Q(\core.CPU_Dmem_value_a5[5][13] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][14]$_SDFFE_PP0P_  (.D(_00565_),
    .Q(\core.CPU_Dmem_value_a5[5][14] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][15]$_SDFFE_PP0P_  (.D(_00566_),
    .Q(\core.CPU_Dmem_value_a5[5][15] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][16]$_SDFFE_PP0P_  (.D(_00567_),
    .Q(\core.CPU_Dmem_value_a5[5][16] ),
    .CLK(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][17]$_SDFFE_PP0P_  (.D(_00568_),
    .Q(\core.CPU_Dmem_value_a5[5][17] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][18]$_SDFFE_PP0P_  (.D(_00569_),
    .Q(\core.CPU_Dmem_value_a5[5][18] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][19]$_SDFFE_PP0P_  (.D(_00570_),
    .Q(\core.CPU_Dmem_value_a5[5][19] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][1]$_SDFFE_PP0P_  (.D(_00571_),
    .Q(\core.CPU_Dmem_value_a5[5][1] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][20]$_SDFFE_PP0P_  (.D(_00572_),
    .Q(\core.CPU_Dmem_value_a5[5][20] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][21]$_SDFFE_PP0P_  (.D(_00573_),
    .Q(\core.CPU_Dmem_value_a5[5][21] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][22]$_SDFFE_PP0P_  (.D(_00574_),
    .Q(\core.CPU_Dmem_value_a5[5][22] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][23]$_SDFFE_PP0P_  (.D(_00575_),
    .Q(\core.CPU_Dmem_value_a5[5][23] ),
    .CLK(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][24]$_SDFFE_PP0P_  (.D(_00576_),
    .Q(\core.CPU_Dmem_value_a5[5][24] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][25]$_SDFFE_PP0P_  (.D(_00577_),
    .Q(\core.CPU_Dmem_value_a5[5][25] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][26]$_SDFFE_PP0P_  (.D(_00578_),
    .Q(\core.CPU_Dmem_value_a5[5][26] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][27]$_SDFFE_PP0P_  (.D(_00579_),
    .Q(\core.CPU_Dmem_value_a5[5][27] ),
    .CLK(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][28]$_SDFFE_PP0P_  (.D(_00580_),
    .Q(\core.CPU_Dmem_value_a5[5][28] ),
    .CLK(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][29]$_SDFFE_PP0P_  (.D(_00581_),
    .Q(\core.CPU_Dmem_value_a5[5][29] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][2]$_SDFFE_PP1P_  (.D(_00582_),
    .Q(\core.CPU_Dmem_value_a5[5][2] ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][30]$_SDFFE_PP0P_  (.D(_00583_),
    .Q(\core.CPU_Dmem_value_a5[5][30] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][31]$_SDFFE_PP0P_  (.D(_00584_),
    .Q(\core.CPU_Dmem_value_a5[5][31] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][3]$_SDFFE_PP0P_  (.D(_00585_),
    .Q(\core.CPU_Dmem_value_a5[5][3] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][4]$_SDFFE_PP0P_  (.D(_00586_),
    .Q(\core.CPU_Dmem_value_a5[5][4] ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][5]$_SDFFE_PP0P_  (.D(_00587_),
    .Q(\core.CPU_Dmem_value_a5[5][5] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][6]$_SDFFE_PP0P_  (.D(_00588_),
    .Q(\core.CPU_Dmem_value_a5[5][6] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][7]$_SDFFE_PP0P_  (.D(_00589_),
    .Q(\core.CPU_Dmem_value_a5[5][7] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][8]$_SDFFE_PP0P_  (.D(_00590_),
    .Q(\core.CPU_Dmem_value_a5[5][8] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[5][9]$_SDFFE_PP0P_  (.D(_00591_),
    .Q(\core.CPU_Dmem_value_a5[5][9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][0]$_SDFFE_PP0P_  (.D(_00592_),
    .Q(\core.CPU_Dmem_value_a5[6][0] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][10]$_SDFFE_PP0P_  (.D(_00593_),
    .Q(\core.CPU_Dmem_value_a5[6][10] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][11]$_SDFFE_PP0P_  (.D(_00594_),
    .Q(\core.CPU_Dmem_value_a5[6][11] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][12]$_SDFFE_PP0P_  (.D(_00595_),
    .Q(\core.CPU_Dmem_value_a5[6][12] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][13]$_SDFFE_PP0P_  (.D(_00596_),
    .Q(\core.CPU_Dmem_value_a5[6][13] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][14]$_SDFFE_PP0P_  (.D(_00597_),
    .Q(\core.CPU_Dmem_value_a5[6][14] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][15]$_SDFFE_PP0P_  (.D(_00598_),
    .Q(\core.CPU_Dmem_value_a5[6][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][16]$_SDFFE_PP0P_  (.D(_00599_),
    .Q(\core.CPU_Dmem_value_a5[6][16] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][17]$_SDFFE_PP0P_  (.D(_00600_),
    .Q(\core.CPU_Dmem_value_a5[6][17] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][18]$_SDFFE_PP0P_  (.D(_00601_),
    .Q(\core.CPU_Dmem_value_a5[6][18] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][19]$_SDFFE_PP0P_  (.D(_00602_),
    .Q(\core.CPU_Dmem_value_a5[6][19] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][1]$_SDFFE_PP1P_  (.D(_00603_),
    .Q(\core.CPU_Dmem_value_a5[6][1] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][20]$_SDFFE_PP0P_  (.D(_00604_),
    .Q(\core.CPU_Dmem_value_a5[6][20] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][21]$_SDFFE_PP0P_  (.D(_00605_),
    .Q(\core.CPU_Dmem_value_a5[6][21] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][22]$_SDFFE_PP0P_  (.D(_00606_),
    .Q(\core.CPU_Dmem_value_a5[6][22] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][23]$_SDFFE_PP0P_  (.D(_00607_),
    .Q(\core.CPU_Dmem_value_a5[6][23] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][24]$_SDFFE_PP0P_  (.D(_00608_),
    .Q(\core.CPU_Dmem_value_a5[6][24] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][25]$_SDFFE_PP0P_  (.D(_00609_),
    .Q(\core.CPU_Dmem_value_a5[6][25] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][26]$_SDFFE_PP0P_  (.D(_00610_),
    .Q(\core.CPU_Dmem_value_a5[6][26] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][27]$_SDFFE_PP0P_  (.D(_00611_),
    .Q(\core.CPU_Dmem_value_a5[6][27] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][28]$_SDFFE_PP0P_  (.D(_00612_),
    .Q(\core.CPU_Dmem_value_a5[6][28] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][29]$_SDFFE_PP0P_  (.D(_00613_),
    .Q(\core.CPU_Dmem_value_a5[6][29] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][2]$_SDFFE_PP1P_  (.D(_00614_),
    .Q(\core.CPU_Dmem_value_a5[6][2] ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][30]$_SDFFE_PP0P_  (.D(_00615_),
    .Q(\core.CPU_Dmem_value_a5[6][30] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][31]$_SDFFE_PP0P_  (.D(_00616_),
    .Q(\core.CPU_Dmem_value_a5[6][31] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][3]$_SDFFE_PP0P_  (.D(_00617_),
    .Q(\core.CPU_Dmem_value_a5[6][3] ),
    .CLK(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][4]$_SDFFE_PP0P_  (.D(_00618_),
    .Q(\core.CPU_Dmem_value_a5[6][4] ),
    .CLK(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][5]$_SDFFE_PP0P_  (.D(_00619_),
    .Q(\core.CPU_Dmem_value_a5[6][5] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][6]$_SDFFE_PP0P_  (.D(_00620_),
    .Q(\core.CPU_Dmem_value_a5[6][6] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][7]$_SDFFE_PP0P_  (.D(_00621_),
    .Q(\core.CPU_Dmem_value_a5[6][7] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][8]$_SDFFE_PP0P_  (.D(_00622_),
    .Q(\core.CPU_Dmem_value_a5[6][8] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[6][9]$_SDFFE_PP0P_  (.D(_00623_),
    .Q(\core.CPU_Dmem_value_a5[6][9] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][0]$_SDFFE_PP1P_  (.D(_00624_),
    .Q(\core.CPU_Dmem_value_a5[7][0] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][10]$_SDFFE_PP0P_  (.D(_00625_),
    .Q(\core.CPU_Dmem_value_a5[7][10] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][11]$_SDFFE_PP0P_  (.D(_00626_),
    .Q(\core.CPU_Dmem_value_a5[7][11] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][12]$_SDFFE_PP0P_  (.D(_00627_),
    .Q(\core.CPU_Dmem_value_a5[7][12] ),
    .CLK(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][13]$_SDFFE_PP0P_  (.D(_00628_),
    .Q(\core.CPU_Dmem_value_a5[7][13] ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][14]$_SDFFE_PP0P_  (.D(_00629_),
    .Q(\core.CPU_Dmem_value_a5[7][14] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][15]$_SDFFE_PP0P_  (.D(_00630_),
    .Q(\core.CPU_Dmem_value_a5[7][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][16]$_SDFFE_PP0P_  (.D(_00631_),
    .Q(\core.CPU_Dmem_value_a5[7][16] ),
    .CLK(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][17]$_SDFFE_PP0P_  (.D(_00632_),
    .Q(\core.CPU_Dmem_value_a5[7][17] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][18]$_SDFFE_PP0P_  (.D(_00633_),
    .Q(\core.CPU_Dmem_value_a5[7][18] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][19]$_SDFFE_PP0P_  (.D(_00634_),
    .Q(\core.CPU_Dmem_value_a5[7][19] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][1]$_SDFFE_PP1P_  (.D(_00635_),
    .Q(\core.CPU_Dmem_value_a5[7][1] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][20]$_SDFFE_PP0P_  (.D(_00636_),
    .Q(\core.CPU_Dmem_value_a5[7][20] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][21]$_SDFFE_PP0P_  (.D(_00637_),
    .Q(\core.CPU_Dmem_value_a5[7][21] ),
    .CLK(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][22]$_SDFFE_PP0P_  (.D(_00638_),
    .Q(\core.CPU_Dmem_value_a5[7][22] ),
    .CLK(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][23]$_SDFFE_PP0P_  (.D(_00639_),
    .Q(\core.CPU_Dmem_value_a5[7][23] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][24]$_SDFFE_PP0P_  (.D(_00640_),
    .Q(\core.CPU_Dmem_value_a5[7][24] ),
    .CLK(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][25]$_SDFFE_PP0P_  (.D(_00641_),
    .Q(\core.CPU_Dmem_value_a5[7][25] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][26]$_SDFFE_PP0P_  (.D(_00642_),
    .Q(\core.CPU_Dmem_value_a5[7][26] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][27]$_SDFFE_PP0P_  (.D(_00643_),
    .Q(\core.CPU_Dmem_value_a5[7][27] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][28]$_SDFFE_PP0P_  (.D(_00644_),
    .Q(\core.CPU_Dmem_value_a5[7][28] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][29]$_SDFFE_PP0P_  (.D(_00645_),
    .Q(\core.CPU_Dmem_value_a5[7][29] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][2]$_SDFFE_PP1P_  (.D(_00646_),
    .Q(\core.CPU_Dmem_value_a5[7][2] ),
    .CLK(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][30]$_SDFFE_PP0P_  (.D(_00647_),
    .Q(\core.CPU_Dmem_value_a5[7][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][31]$_SDFFE_PP0P_  (.D(_00648_),
    .Q(\core.CPU_Dmem_value_a5[7][31] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][3]$_SDFFE_PP0P_  (.D(_00649_),
    .Q(\core.CPU_Dmem_value_a5[7][3] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][4]$_SDFFE_PP0P_  (.D(_00650_),
    .Q(\core.CPU_Dmem_value_a5[7][4] ),
    .CLK(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][5]$_SDFFE_PP0P_  (.D(_00651_),
    .Q(\core.CPU_Dmem_value_a5[7][5] ),
    .CLK(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][6]$_SDFFE_PP0P_  (.D(_00652_),
    .Q(\core.CPU_Dmem_value_a5[7][6] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][7]$_SDFFE_PP0P_  (.D(_00653_),
    .Q(\core.CPU_Dmem_value_a5[7][7] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][8]$_SDFFE_PP0P_  (.D(_00654_),
    .Q(\core.CPU_Dmem_value_a5[7][8] ),
    .CLK(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[7][9]$_SDFFE_PP0P_  (.D(_00655_),
    .Q(\core.CPU_Dmem_value_a5[7][9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][0]$_SDFFE_PP0P_  (.D(_00656_),
    .Q(\core.CPU_Dmem_value_a5[8][0] ),
    .CLK(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][10]$_SDFFE_PP0P_  (.D(_00657_),
    .Q(\core.CPU_Dmem_value_a5[8][10] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][11]$_SDFFE_PP0P_  (.D(_00658_),
    .Q(\core.CPU_Dmem_value_a5[8][11] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][12]$_SDFFE_PP0P_  (.D(_00659_),
    .Q(\core.CPU_Dmem_value_a5[8][12] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][13]$_SDFFE_PP0P_  (.D(_00660_),
    .Q(\core.CPU_Dmem_value_a5[8][13] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][14]$_SDFFE_PP0P_  (.D(_00661_),
    .Q(\core.CPU_Dmem_value_a5[8][14] ),
    .CLK(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][15]$_SDFFE_PP0P_  (.D(_00662_),
    .Q(\core.CPU_Dmem_value_a5[8][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][16]$_SDFFE_PP0P_  (.D(_00663_),
    .Q(\core.CPU_Dmem_value_a5[8][16] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][17]$_SDFFE_PP0P_  (.D(_00664_),
    .Q(\core.CPU_Dmem_value_a5[8][17] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][18]$_SDFFE_PP0P_  (.D(_00665_),
    .Q(\core.CPU_Dmem_value_a5[8][18] ),
    .CLK(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][19]$_SDFFE_PP0P_  (.D(_00666_),
    .Q(\core.CPU_Dmem_value_a5[8][19] ),
    .CLK(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][1]$_SDFFE_PP0P_  (.D(_00667_),
    .Q(\core.CPU_Dmem_value_a5[8][1] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][20]$_SDFFE_PP0P_  (.D(_00668_),
    .Q(\core.CPU_Dmem_value_a5[8][20] ),
    .CLK(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][21]$_SDFFE_PP0P_  (.D(_00669_),
    .Q(\core.CPU_Dmem_value_a5[8][21] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][22]$_SDFFE_PP0P_  (.D(_00670_),
    .Q(\core.CPU_Dmem_value_a5[8][22] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][23]$_SDFFE_PP0P_  (.D(_00671_),
    .Q(\core.CPU_Dmem_value_a5[8][23] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][24]$_SDFFE_PP0P_  (.D(_00672_),
    .Q(\core.CPU_Dmem_value_a5[8][24] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][25]$_SDFFE_PP0P_  (.D(_00673_),
    .Q(\core.CPU_Dmem_value_a5[8][25] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][26]$_SDFFE_PP0P_  (.D(_00674_),
    .Q(\core.CPU_Dmem_value_a5[8][26] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][27]$_SDFFE_PP0P_  (.D(_00675_),
    .Q(\core.CPU_Dmem_value_a5[8][27] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][28]$_SDFFE_PP0P_  (.D(_00676_),
    .Q(\core.CPU_Dmem_value_a5[8][28] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][29]$_SDFFE_PP0P_  (.D(_00677_),
    .Q(\core.CPU_Dmem_value_a5[8][29] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][2]$_SDFFE_PP0P_  (.D(_00678_),
    .Q(\core.CPU_Dmem_value_a5[8][2] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][30]$_SDFFE_PP0P_  (.D(_00679_),
    .Q(\core.CPU_Dmem_value_a5[8][30] ),
    .CLK(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][31]$_SDFFE_PP0P_  (.D(_00680_),
    .Q(\core.CPU_Dmem_value_a5[8][31] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][3]$_SDFFE_PP1P_  (.D(_00681_),
    .Q(\core.CPU_Dmem_value_a5[8][3] ),
    .CLK(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][4]$_SDFFE_PP0P_  (.D(_00682_),
    .Q(\core.CPU_Dmem_value_a5[8][4] ),
    .CLK(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][5]$_SDFFE_PP0P_  (.D(_00683_),
    .Q(\core.CPU_Dmem_value_a5[8][5] ),
    .CLK(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][6]$_SDFFE_PP0P_  (.D(_00684_),
    .Q(\core.CPU_Dmem_value_a5[8][6] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][7]$_SDFFE_PP0P_  (.D(_00685_),
    .Q(\core.CPU_Dmem_value_a5[8][7] ),
    .CLK(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][8]$_SDFFE_PP0P_  (.D(_00686_),
    .Q(\core.CPU_Dmem_value_a5[8][8] ),
    .CLK(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[8][9]$_SDFFE_PP0P_  (.D(_00687_),
    .Q(\core.CPU_Dmem_value_a5[8][9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][0]$_SDFFE_PP1P_  (.D(_00688_),
    .Q(\core.CPU_Dmem_value_a5[9][0] ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][10]$_SDFFE_PP0P_  (.D(_00689_),
    .Q(\core.CPU_Dmem_value_a5[9][10] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][11]$_SDFFE_PP0P_  (.D(_00690_),
    .Q(\core.CPU_Dmem_value_a5[9][11] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][12]$_SDFFE_PP0P_  (.D(_00691_),
    .Q(\core.CPU_Dmem_value_a5[9][12] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][13]$_SDFFE_PP0P_  (.D(_00692_),
    .Q(\core.CPU_Dmem_value_a5[9][13] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][14]$_SDFFE_PP0P_  (.D(_00693_),
    .Q(\core.CPU_Dmem_value_a5[9][14] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][15]$_SDFFE_PP0P_  (.D(_00694_),
    .Q(\core.CPU_Dmem_value_a5[9][15] ),
    .CLK(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][16]$_SDFFE_PP0P_  (.D(_00695_),
    .Q(\core.CPU_Dmem_value_a5[9][16] ),
    .CLK(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][17]$_SDFFE_PP0P_  (.D(_00696_),
    .Q(\core.CPU_Dmem_value_a5[9][17] ),
    .CLK(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][18]$_SDFFE_PP0P_  (.D(_00697_),
    .Q(\core.CPU_Dmem_value_a5[9][18] ),
    .CLK(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][19]$_SDFFE_PP0P_  (.D(_00698_),
    .Q(\core.CPU_Dmem_value_a5[9][19] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][1]$_SDFFE_PP0P_  (.D(_00699_),
    .Q(\core.CPU_Dmem_value_a5[9][1] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][20]$_SDFFE_PP0P_  (.D(_00700_),
    .Q(\core.CPU_Dmem_value_a5[9][20] ),
    .CLK(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][21]$_SDFFE_PP0P_  (.D(_00701_),
    .Q(\core.CPU_Dmem_value_a5[9][21] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][22]$_SDFFE_PP0P_  (.D(_00702_),
    .Q(\core.CPU_Dmem_value_a5[9][22] ),
    .CLK(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][23]$_SDFFE_PP0P_  (.D(_00703_),
    .Q(\core.CPU_Dmem_value_a5[9][23] ),
    .CLK(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][24]$_SDFFE_PP0P_  (.D(_00704_),
    .Q(\core.CPU_Dmem_value_a5[9][24] ),
    .CLK(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][25]$_SDFFE_PP0P_  (.D(_00705_),
    .Q(\core.CPU_Dmem_value_a5[9][25] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][26]$_SDFFE_PP0P_  (.D(_00706_),
    .Q(\core.CPU_Dmem_value_a5[9][26] ),
    .CLK(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][27]$_SDFFE_PP0P_  (.D(_00707_),
    .Q(\core.CPU_Dmem_value_a5[9][27] ),
    .CLK(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][28]$_SDFFE_PP0P_  (.D(_00708_),
    .Q(\core.CPU_Dmem_value_a5[9][28] ),
    .CLK(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][29]$_SDFFE_PP0P_  (.D(_00709_),
    .Q(\core.CPU_Dmem_value_a5[9][29] ),
    .CLK(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][2]$_SDFFE_PP0P_  (.D(_00710_),
    .Q(\core.CPU_Dmem_value_a5[9][2] ),
    .CLK(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][30]$_SDFFE_PP0P_  (.D(_00711_),
    .Q(\core.CPU_Dmem_value_a5[9][30] ),
    .CLK(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][31]$_SDFFE_PP0P_  (.D(_00712_),
    .Q(\core.CPU_Dmem_value_a5[9][31] ),
    .CLK(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][3]$_SDFFE_PP1P_  (.D(_00713_),
    .Q(\core.CPU_Dmem_value_a5[9][3] ),
    .CLK(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][4]$_SDFFE_PP0P_  (.D(_00714_),
    .Q(\core.CPU_Dmem_value_a5[9][4] ),
    .CLK(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][5]$_SDFFE_PP0P_  (.D(_00715_),
    .Q(\core.CPU_Dmem_value_a5[9][5] ),
    .CLK(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][6]$_SDFFE_PP0P_  (.D(_00716_),
    .Q(\core.CPU_Dmem_value_a5[9][6] ),
    .CLK(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][7]$_SDFFE_PP0P_  (.D(_00717_),
    .Q(\core.CPU_Dmem_value_a5[9][7] ),
    .CLK(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][8]$_SDFFE_PP0P_  (.D(_00718_),
    .Q(\core.CPU_Dmem_value_a5[9][8] ),
    .CLK(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Dmem_value_a5[9][9]$_SDFFE_PP0P_  (.D(_00719_),
    .Q(\core.CPU_Dmem_value_a5[9][9] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][0]$_SDFFE_PP0P_  (.D(_00720_),
    .Q(\core.CPU_Xreg_value_a4[0][0] ),
    .CLK(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][10]$_SDFFE_PP0P_  (.D(_00721_),
    .Q(\core.CPU_Xreg_value_a4[0][10] ),
    .CLK(clknet_leaf_110_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][11]$_SDFFE_PP0P_  (.D(_00722_),
    .Q(\core.CPU_Xreg_value_a4[0][11] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][12]$_SDFFE_PP0P_  (.D(_00723_),
    .Q(\core.CPU_Xreg_value_a4[0][12] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][13]$_SDFFE_PP0P_  (.D(_00724_),
    .Q(\core.CPU_Xreg_value_a4[0][13] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][14]$_SDFFE_PP0P_  (.D(_00725_),
    .Q(\core.CPU_Xreg_value_a4[0][14] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][15]$_SDFFE_PP0P_  (.D(_00726_),
    .Q(\core.CPU_Xreg_value_a4[0][15] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][16]$_SDFFE_PP0P_  (.D(_00727_),
    .Q(\core.CPU_Xreg_value_a4[0][16] ),
    .CLK(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][17]$_SDFFE_PP0P_  (.D(_00728_),
    .Q(\core.CPU_Xreg_value_a4[0][17] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][18]$_SDFFE_PP0P_  (.D(_00729_),
    .Q(\core.CPU_Xreg_value_a4[0][18] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][19]$_SDFFE_PP0P_  (.D(_00730_),
    .Q(\core.CPU_Xreg_value_a4[0][19] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][1]$_SDFFE_PP0P_  (.D(_00731_),
    .Q(\core.CPU_Xreg_value_a4[0][1] ),
    .CLK(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][20]$_SDFFE_PP0P_  (.D(_00732_),
    .Q(\core.CPU_Xreg_value_a4[0][20] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][21]$_SDFFE_PP0P_  (.D(_00733_),
    .Q(\core.CPU_Xreg_value_a4[0][21] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][22]$_SDFFE_PP0P_  (.D(_00734_),
    .Q(\core.CPU_Xreg_value_a4[0][22] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][23]$_SDFFE_PP0P_  (.D(_00735_),
    .Q(\core.CPU_Xreg_value_a4[0][23] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][24]$_SDFFE_PP0P_  (.D(_00736_),
    .Q(\core.CPU_Xreg_value_a4[0][24] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][25]$_SDFFE_PP0P_  (.D(_00737_),
    .Q(\core.CPU_Xreg_value_a4[0][25] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][26]$_SDFFE_PP0P_  (.D(_00738_),
    .Q(\core.CPU_Xreg_value_a4[0][26] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][27]$_SDFFE_PP0P_  (.D(_00739_),
    .Q(\core.CPU_Xreg_value_a4[0][27] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][28]$_SDFFE_PP0P_  (.D(_00740_),
    .Q(\core.CPU_Xreg_value_a4[0][28] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][29]$_SDFFE_PP0P_  (.D(_00741_),
    .Q(\core.CPU_Xreg_value_a4[0][29] ),
    .CLK(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][2]$_SDFFE_PP0P_  (.D(_00742_),
    .Q(\core.CPU_Xreg_value_a4[0][2] ),
    .CLK(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][30]$_SDFFE_PP0P_  (.D(_00743_),
    .Q(\core.CPU_Xreg_value_a4[0][30] ),
    .CLK(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][31]$_SDFFE_PP0P_  (.D(_00744_),
    .Q(\core.CPU_Xreg_value_a4[0][31] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][3]$_SDFFE_PP0P_  (.D(_00745_),
    .Q(\core.CPU_Xreg_value_a4[0][3] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][4]$_SDFFE_PP0P_  (.D(_00746_),
    .Q(\core.CPU_Xreg_value_a4[0][4] ),
    .CLK(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][5]$_SDFFE_PP0P_  (.D(_00747_),
    .Q(\core.CPU_Xreg_value_a4[0][5] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][6]$_SDFFE_PP0P_  (.D(_00748_),
    .Q(\core.CPU_Xreg_value_a4[0][6] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][7]$_SDFFE_PP0P_  (.D(_00749_),
    .Q(\core.CPU_Xreg_value_a4[0][7] ),
    .CLK(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][8]$_SDFFE_PP0P_  (.D(_00750_),
    .Q(\core.CPU_Xreg_value_a4[0][8] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[0][9]$_SDFFE_PP0P_  (.D(_00751_),
    .Q(\core.CPU_Xreg_value_a4[0][9] ),
    .CLK(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][0]$_SDFFE_PP0P_  (.D(_00752_),
    .Q(\core.CPU_Xreg_value_a4[10][0] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][10]$_SDFFE_PP0P_  (.D(_00753_),
    .Q(\core.CPU_Xreg_value_a4[10][10] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][11]$_SDFFE_PP0P_  (.D(_00754_),
    .Q(\core.CPU_Xreg_value_a4[10][11] ),
    .CLK(clknet_leaf_110_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][12]$_SDFFE_PP0P_  (.D(_00755_),
    .Q(\core.CPU_Xreg_value_a4[10][12] ),
    .CLK(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][13]$_SDFFE_PP0P_  (.D(_00756_),
    .Q(\core.CPU_Xreg_value_a4[10][13] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][14]$_SDFFE_PP0P_  (.D(_00757_),
    .Q(\core.CPU_Xreg_value_a4[10][14] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][15]$_SDFFE_PP0P_  (.D(_00758_),
    .Q(\core.CPU_Xreg_value_a4[10][15] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][16]$_SDFFE_PP0P_  (.D(_00759_),
    .Q(\core.CPU_Xreg_value_a4[10][16] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][17]$_SDFFE_PP0P_  (.D(_00760_),
    .Q(\core.CPU_Xreg_value_a4[10][17] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][18]$_SDFFE_PP0P_  (.D(_00761_),
    .Q(\core.CPU_Xreg_value_a4[10][18] ),
    .CLK(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][19]$_SDFFE_PP0P_  (.D(_00762_),
    .Q(\core.CPU_Xreg_value_a4[10][19] ),
    .CLK(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][1]$_SDFFE_PP1P_  (.D(_00763_),
    .Q(\core.CPU_Xreg_value_a4[10][1] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][20]$_SDFFE_PP0P_  (.D(_00764_),
    .Q(\core.CPU_Xreg_value_a4[10][20] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][21]$_SDFFE_PP0P_  (.D(_00765_),
    .Q(\core.CPU_Xreg_value_a4[10][21] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][22]$_SDFFE_PP0P_  (.D(_00766_),
    .Q(\core.CPU_Xreg_value_a4[10][22] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][23]$_SDFFE_PP0P_  (.D(_00767_),
    .Q(\core.CPU_Xreg_value_a4[10][23] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][24]$_SDFFE_PP0P_  (.D(_00768_),
    .Q(\core.CPU_Xreg_value_a4[10][24] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][25]$_SDFFE_PP0P_  (.D(_00769_),
    .Q(\core.CPU_Xreg_value_a4[10][25] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][26]$_SDFFE_PP0P_  (.D(_00770_),
    .Q(\core.CPU_Xreg_value_a4[10][26] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][27]$_SDFFE_PP0P_  (.D(_00771_),
    .Q(\core.CPU_Xreg_value_a4[10][27] ),
    .CLK(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][28]$_SDFFE_PP0P_  (.D(_00772_),
    .Q(\core.CPU_Xreg_value_a4[10][28] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][29]$_SDFFE_PP0P_  (.D(_00773_),
    .Q(\core.CPU_Xreg_value_a4[10][29] ),
    .CLK(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][2]$_SDFFE_PP0P_  (.D(_00774_),
    .Q(\core.CPU_Xreg_value_a4[10][2] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][30]$_SDFFE_PP0P_  (.D(_00775_),
    .Q(\core.CPU_Xreg_value_a4[10][30] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][31]$_SDFFE_PP0P_  (.D(_00776_),
    .Q(\core.CPU_Xreg_value_a4[10][31] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][3]$_SDFFE_PP1P_  (.D(_00777_),
    .Q(\core.CPU_Xreg_value_a4[10][3] ),
    .CLK(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][4]$_SDFFE_PP0P_  (.D(_00778_),
    .Q(\core.CPU_Xreg_value_a4[10][4] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][5]$_SDFFE_PP0P_  (.D(_00779_),
    .Q(\core.CPU_Xreg_value_a4[10][5] ),
    .CLK(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][6]$_SDFFE_PP0P_  (.D(_00780_),
    .Q(\core.CPU_Xreg_value_a4[10][6] ),
    .CLK(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][7]$_SDFFE_PP0P_  (.D(_00781_),
    .Q(\core.CPU_Xreg_value_a4[10][7] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][8]$_SDFFE_PP0P_  (.D(_00782_),
    .Q(\core.CPU_Xreg_value_a4[10][8] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[10][9]$_SDFFE_PP0P_  (.D(_00783_),
    .Q(\core.CPU_Xreg_value_a4[10][9] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][0]$_SDFFE_PP1P_  (.D(_00784_),
    .Q(\core.CPU_Xreg_value_a4[11][0] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][10]$_SDFFE_PP0P_  (.D(_00785_),
    .Q(\core.CPU_Xreg_value_a4[11][10] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][11]$_SDFFE_PP0P_  (.D(_00786_),
    .Q(\core.CPU_Xreg_value_a4[11][11] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][12]$_SDFFE_PP0P_  (.D(_00787_),
    .Q(\core.CPU_Xreg_value_a4[11][12] ),
    .CLK(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][13]$_SDFFE_PP0P_  (.D(_00788_),
    .Q(\core.CPU_Xreg_value_a4[11][13] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][14]$_SDFFE_PP0P_  (.D(_00789_),
    .Q(\core.CPU_Xreg_value_a4[11][14] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][15]$_SDFFE_PP0P_  (.D(_00790_),
    .Q(\core.CPU_Xreg_value_a4[11][15] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][16]$_SDFFE_PP0P_  (.D(_00791_),
    .Q(\core.CPU_Xreg_value_a4[11][16] ),
    .CLK(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][17]$_SDFFE_PP0P_  (.D(_00792_),
    .Q(\core.CPU_Xreg_value_a4[11][17] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][18]$_SDFFE_PP0P_  (.D(_00793_),
    .Q(\core.CPU_Xreg_value_a4[11][18] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][19]$_SDFFE_PP0P_  (.D(_00794_),
    .Q(\core.CPU_Xreg_value_a4[11][19] ),
    .CLK(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][1]$_SDFFE_PP1P_  (.D(_00795_),
    .Q(\core.CPU_Xreg_value_a4[11][1] ),
    .CLK(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][20]$_SDFFE_PP0P_  (.D(_00796_),
    .Q(\core.CPU_Xreg_value_a4[11][20] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][21]$_SDFFE_PP0P_  (.D(_00797_),
    .Q(\core.CPU_Xreg_value_a4[11][21] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][22]$_SDFFE_PP0P_  (.D(_00798_),
    .Q(\core.CPU_Xreg_value_a4[11][22] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][23]$_SDFFE_PP0P_  (.D(_00799_),
    .Q(\core.CPU_Xreg_value_a4[11][23] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][24]$_SDFFE_PP0P_  (.D(_00800_),
    .Q(\core.CPU_Xreg_value_a4[11][24] ),
    .CLK(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][25]$_SDFFE_PP0P_  (.D(_00801_),
    .Q(\core.CPU_Xreg_value_a4[11][25] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][26]$_SDFFE_PP0P_  (.D(_00802_),
    .Q(\core.CPU_Xreg_value_a4[11][26] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][27]$_SDFFE_PP0P_  (.D(_00803_),
    .Q(\core.CPU_Xreg_value_a4[11][27] ),
    .CLK(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][28]$_SDFFE_PP0P_  (.D(_00804_),
    .Q(\core.CPU_Xreg_value_a4[11][28] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][29]$_SDFFE_PP0P_  (.D(_00805_),
    .Q(\core.CPU_Xreg_value_a4[11][29] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][2]$_SDFFE_PP0P_  (.D(_00806_),
    .Q(\core.CPU_Xreg_value_a4[11][2] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][30]$_SDFFE_PP0P_  (.D(_00807_),
    .Q(\core.CPU_Xreg_value_a4[11][30] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][31]$_SDFFE_PP0P_  (.D(_00808_),
    .Q(\core.CPU_Xreg_value_a4[11][31] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][3]$_SDFFE_PP1P_  (.D(_00809_),
    .Q(\core.CPU_Xreg_value_a4[11][3] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][4]$_SDFFE_PP0P_  (.D(_00810_),
    .Q(\core.CPU_Xreg_value_a4[11][4] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][5]$_SDFFE_PP0P_  (.D(_00811_),
    .Q(\core.CPU_Xreg_value_a4[11][5] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][6]$_SDFFE_PP0P_  (.D(_00812_),
    .Q(\core.CPU_Xreg_value_a4[11][6] ),
    .CLK(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][7]$_SDFFE_PP0P_  (.D(_00813_),
    .Q(\core.CPU_Xreg_value_a4[11][7] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][8]$_SDFFE_PP0P_  (.D(_00814_),
    .Q(\core.CPU_Xreg_value_a4[11][8] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[11][9]$_SDFFE_PP0P_  (.D(_00815_),
    .Q(\core.CPU_Xreg_value_a4[11][9] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][0]$_SDFFE_PP0P_  (.D(_00816_),
    .Q(\core.CPU_Xreg_value_a4[16][0] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][10]$_SDFFE_PP0P_  (.D(_00817_),
    .Q(\core.CPU_Xreg_value_a4[16][10] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][11]$_SDFFE_PP0P_  (.D(_00818_),
    .Q(\core.CPU_Xreg_value_a4[16][11] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][12]$_SDFFE_PP0P_  (.D(_00819_),
    .Q(\core.CPU_Xreg_value_a4[16][12] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][13]$_SDFFE_PP0P_  (.D(_00820_),
    .Q(\core.CPU_Xreg_value_a4[16][13] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][14]$_SDFFE_PP0P_  (.D(_00821_),
    .Q(\core.CPU_Xreg_value_a4[16][14] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][15]$_SDFFE_PP0P_  (.D(_00822_),
    .Q(\core.CPU_Xreg_value_a4[16][15] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][16]$_SDFFE_PP0P_  (.D(_00823_),
    .Q(\core.CPU_Xreg_value_a4[16][16] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][17]$_SDFFE_PP0P_  (.D(_00824_),
    .Q(\core.CPU_Xreg_value_a4[16][17] ),
    .CLK(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][18]$_SDFFE_PP0P_  (.D(_00825_),
    .Q(\core.CPU_Xreg_value_a4[16][18] ),
    .CLK(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][19]$_SDFFE_PP0P_  (.D(_00826_),
    .Q(\core.CPU_Xreg_value_a4[16][19] ),
    .CLK(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][1]$_SDFFE_PP0P_  (.D(_00827_),
    .Q(\core.CPU_Xreg_value_a4[16][1] ),
    .CLK(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][20]$_SDFFE_PP0P_  (.D(_00828_),
    .Q(\core.CPU_Xreg_value_a4[16][20] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][21]$_SDFFE_PP0P_  (.D(_00829_),
    .Q(\core.CPU_Xreg_value_a4[16][21] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][22]$_SDFFE_PP0P_  (.D(_00830_),
    .Q(\core.CPU_Xreg_value_a4[16][22] ),
    .CLK(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][23]$_SDFFE_PP0P_  (.D(_00831_),
    .Q(\core.CPU_Xreg_value_a4[16][23] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][24]$_SDFFE_PP0P_  (.D(_00832_),
    .Q(\core.CPU_Xreg_value_a4[16][24] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][25]$_SDFFE_PP0P_  (.D(_00833_),
    .Q(\core.CPU_Xreg_value_a4[16][25] ),
    .CLK(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][26]$_SDFFE_PP0P_  (.D(_00834_),
    .Q(\core.CPU_Xreg_value_a4[16][26] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][27]$_SDFFE_PP0P_  (.D(_00835_),
    .Q(\core.CPU_Xreg_value_a4[16][27] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][28]$_SDFFE_PP0P_  (.D(_00836_),
    .Q(\core.CPU_Xreg_value_a4[16][28] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][29]$_SDFFE_PP0P_  (.D(_00837_),
    .Q(\core.CPU_Xreg_value_a4[16][29] ),
    .CLK(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][2]$_SDFFE_PP0P_  (.D(_00838_),
    .Q(\core.CPU_Xreg_value_a4[16][2] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][30]$_SDFFE_PP0P_  (.D(_00839_),
    .Q(\core.CPU_Xreg_value_a4[16][30] ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][31]$_SDFFE_PP0P_  (.D(_00840_),
    .Q(\core.CPU_Xreg_value_a4[16][31] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][3]$_SDFFE_PP0P_  (.D(_00841_),
    .Q(\core.CPU_Xreg_value_a4[16][3] ),
    .CLK(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][4]$_SDFFE_PP1P_  (.D(_00842_),
    .Q(\core.CPU_Xreg_value_a4[16][4] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][5]$_SDFFE_PP0P_  (.D(_00843_),
    .Q(\core.CPU_Xreg_value_a4[16][5] ),
    .CLK(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][6]$_SDFFE_PP0P_  (.D(_00844_),
    .Q(\core.CPU_Xreg_value_a4[16][6] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][7]$_SDFFE_PP0P_  (.D(_00845_),
    .Q(\core.CPU_Xreg_value_a4[16][7] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][8]$_SDFFE_PP0P_  (.D(_00846_),
    .Q(\core.CPU_Xreg_value_a4[16][8] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[16][9]$_SDFFE_PP0P_  (.D(_00847_),
    .Q(\core.CPU_Xreg_value_a4[16][9] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][0]$_SDFFE_PP1P_  (.D(_00848_),
    .Q(\core.CPU_Xreg_value_a4[17][0] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][10]$_SDFFE_PP0P_  (.D(_00849_),
    .Q(\core.CPU_Xreg_value_a4[17][10] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][11]$_SDFFE_PP0P_  (.D(_00850_),
    .Q(\core.CPU_Xreg_value_a4[17][11] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][12]$_SDFFE_PP0P_  (.D(_00851_),
    .Q(\core.CPU_Xreg_value_a4[17][12] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][13]$_SDFFE_PP0P_  (.D(_00852_),
    .Q(\core.CPU_Xreg_value_a4[17][13] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][14]$_SDFFE_PP0P_  (.D(_00853_),
    .Q(\core.CPU_Xreg_value_a4[17][14] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][15]$_SDFFE_PP0P_  (.D(_00854_),
    .Q(\core.CPU_Xreg_value_a4[17][15] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][16]$_SDFFE_PP0P_  (.D(_00855_),
    .Q(\core.CPU_Xreg_value_a4[17][16] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][17]$_SDFFE_PP0P_  (.D(_00856_),
    .Q(\core.CPU_Xreg_value_a4[17][17] ),
    .CLK(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][18]$_SDFFE_PP0P_  (.D(_00857_),
    .Q(\core.CPU_Xreg_value_a4[17][18] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][19]$_SDFFE_PP0P_  (.D(_00858_),
    .Q(\core.CPU_Xreg_value_a4[17][19] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][1]$_SDFFE_PP0P_  (.D(_00859_),
    .Q(\core.CPU_Xreg_value_a4[17][1] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][20]$_SDFFE_PP0P_  (.D(_00860_),
    .Q(\core.CPU_Xreg_value_a4[17][20] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][21]$_SDFFE_PP0P_  (.D(_00861_),
    .Q(\core.CPU_Xreg_value_a4[17][21] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][22]$_SDFFE_PP0P_  (.D(_00862_),
    .Q(\core.CPU_Xreg_value_a4[17][22] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][23]$_SDFFE_PP0P_  (.D(_00863_),
    .Q(\core.CPU_Xreg_value_a4[17][23] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][24]$_SDFFE_PP0P_  (.D(_00864_),
    .Q(\core.CPU_Xreg_value_a4[17][24] ),
    .CLK(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][25]$_SDFFE_PP0P_  (.D(_00865_),
    .Q(\core.CPU_Xreg_value_a4[17][25] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][26]$_SDFFE_PP0P_  (.D(_00866_),
    .Q(\core.CPU_Xreg_value_a4[17][26] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][27]$_SDFFE_PP0P_  (.D(_00867_),
    .Q(\core.CPU_Xreg_value_a4[17][27] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][28]$_SDFFE_PP0P_  (.D(_00868_),
    .Q(\core.CPU_Xreg_value_a4[17][28] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][29]$_SDFFE_PP0P_  (.D(_00869_),
    .Q(\core.CPU_Xreg_value_a4[17][29] ),
    .CLK(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][2]$_SDFFE_PP0P_  (.D(_00870_),
    .Q(\core.CPU_Xreg_value_a4[17][2] ),
    .CLK(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][30]$_SDFFE_PP0P_  (.D(_00871_),
    .Q(\core.CPU_Xreg_value_a4[17][30] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][31]$_SDFFE_PP0P_  (.D(_00872_),
    .Q(\core.CPU_Xreg_value_a4[17][31] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][3]$_SDFFE_PP0P_  (.D(_00873_),
    .Q(\core.CPU_Xreg_value_a4[17][3] ),
    .CLK(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][4]$_SDFFE_PP1P_  (.D(_00874_),
    .Q(\core.CPU_Xreg_value_a4[17][4] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][5]$_SDFFE_PP0P_  (.D(_00875_),
    .Q(\core.CPU_Xreg_value_a4[17][5] ),
    .CLK(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][6]$_SDFFE_PP0P_  (.D(_00876_),
    .Q(\core.CPU_Xreg_value_a4[17][6] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][7]$_SDFFE_PP0P_  (.D(_00877_),
    .Q(\core.CPU_Xreg_value_a4[17][7] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][8]$_SDFFE_PP0P_  (.D(_00878_),
    .Q(\core.CPU_Xreg_value_a4[17][8] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[17][9]$_SDFFE_PP0P_  (.D(_00879_),
    .Q(\core.CPU_Xreg_value_a4[17][9] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][0]$_SDFFE_PP1P_  (.D(_00880_),
    .Q(\core.CPU_Xreg_value_a4[1][0] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][10]$_SDFFE_PP0P_  (.D(_00881_),
    .Q(\core.CPU_Xreg_value_a4[1][10] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][11]$_SDFFE_PP0P_  (.D(_00882_),
    .Q(\core.CPU_Xreg_value_a4[1][11] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][12]$_SDFFE_PP0P_  (.D(_00883_),
    .Q(\core.CPU_Xreg_value_a4[1][12] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][13]$_SDFFE_PP0P_  (.D(_00884_),
    .Q(\core.CPU_Xreg_value_a4[1][13] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][14]$_SDFFE_PP0P_  (.D(_00885_),
    .Q(\core.CPU_Xreg_value_a4[1][14] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][15]$_SDFFE_PP0P_  (.D(_00886_),
    .Q(\core.CPU_Xreg_value_a4[1][15] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][16]$_SDFFE_PP0P_  (.D(_00887_),
    .Q(\core.CPU_Xreg_value_a4[1][16] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][17]$_SDFFE_PP0P_  (.D(_00888_),
    .Q(\core.CPU_Xreg_value_a4[1][17] ),
    .CLK(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][18]$_SDFFE_PP0P_  (.D(_00889_),
    .Q(\core.CPU_Xreg_value_a4[1][18] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][19]$_SDFFE_PP0P_  (.D(_00890_),
    .Q(\core.CPU_Xreg_value_a4[1][19] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][1]$_SDFFE_PP0P_  (.D(_00891_),
    .Q(\core.CPU_Xreg_value_a4[1][1] ),
    .CLK(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][20]$_SDFFE_PP0P_  (.D(_00892_),
    .Q(\core.CPU_Xreg_value_a4[1][20] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][21]$_SDFFE_PP0P_  (.D(_00893_),
    .Q(\core.CPU_Xreg_value_a4[1][21] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][22]$_SDFFE_PP0P_  (.D(_00894_),
    .Q(\core.CPU_Xreg_value_a4[1][22] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][23]$_SDFFE_PP0P_  (.D(_00895_),
    .Q(\core.CPU_Xreg_value_a4[1][23] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][24]$_SDFFE_PP0P_  (.D(_00896_),
    .Q(\core.CPU_Xreg_value_a4[1][24] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][25]$_SDFFE_PP0P_  (.D(_00897_),
    .Q(\core.CPU_Xreg_value_a4[1][25] ),
    .CLK(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][26]$_SDFFE_PP0P_  (.D(_00898_),
    .Q(\core.CPU_Xreg_value_a4[1][26] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][27]$_SDFFE_PP0P_  (.D(_00899_),
    .Q(\core.CPU_Xreg_value_a4[1][27] ),
    .CLK(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][28]$_SDFFE_PP0P_  (.D(_00900_),
    .Q(\core.CPU_Xreg_value_a4[1][28] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][29]$_SDFFE_PP0P_  (.D(_00901_),
    .Q(\core.CPU_Xreg_value_a4[1][29] ),
    .CLK(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][2]$_SDFFE_PP0P_  (.D(_00902_),
    .Q(\core.CPU_Xreg_value_a4[1][2] ),
    .CLK(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][30]$_SDFFE_PP0P_  (.D(_00903_),
    .Q(\core.CPU_Xreg_value_a4[1][30] ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][31]$_SDFFE_PP0P_  (.D(_00904_),
    .Q(\core.CPU_Xreg_value_a4[1][31] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][3]$_SDFFE_PP0P_  (.D(_00905_),
    .Q(\core.CPU_Xreg_value_a4[1][3] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][4]$_SDFFE_PP0P_  (.D(_00906_),
    .Q(\core.CPU_Xreg_value_a4[1][4] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][5]$_SDFFE_PP0P_  (.D(_00907_),
    .Q(\core.CPU_Xreg_value_a4[1][5] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][6]$_SDFFE_PP0P_  (.D(_00908_),
    .Q(\core.CPU_Xreg_value_a4[1][6] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][7]$_SDFFE_PP0P_  (.D(_00909_),
    .Q(\core.CPU_Xreg_value_a4[1][7] ),
    .CLK(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][8]$_SDFFE_PP0P_  (.D(_00910_),
    .Q(\core.CPU_Xreg_value_a4[1][8] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[1][9]$_SDFFE_PP0P_  (.D(_00911_),
    .Q(\core.CPU_Xreg_value_a4[1][9] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][0]$_SDFFE_PP0P_  (.D(_00912_),
    .Q(\core.CPU_Xreg_value_a4[26][0] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][10]$_SDFFE_PP0P_  (.D(_00913_),
    .Q(\core.CPU_Xreg_value_a4[26][10] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][11]$_SDFFE_PP0P_  (.D(_00914_),
    .Q(\core.CPU_Xreg_value_a4[26][11] ),
    .CLK(clknet_leaf_110_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][12]$_SDFFE_PP0P_  (.D(_00915_),
    .Q(\core.CPU_Xreg_value_a4[26][12] ),
    .CLK(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][13]$_SDFFE_PP0P_  (.D(_00916_),
    .Q(\core.CPU_Xreg_value_a4[26][13] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][14]$_SDFFE_PP0P_  (.D(_00917_),
    .Q(\core.CPU_Xreg_value_a4[26][14] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][15]$_SDFFE_PP0P_  (.D(_00918_),
    .Q(\core.CPU_Xreg_value_a4[26][15] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][16]$_SDFFE_PP0P_  (.D(_00919_),
    .Q(\core.CPU_Xreg_value_a4[26][16] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][17]$_SDFFE_PP0P_  (.D(_00920_),
    .Q(\core.CPU_Xreg_value_a4[26][17] ),
    .CLK(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][18]$_SDFFE_PP0P_  (.D(_00921_),
    .Q(\core.CPU_Xreg_value_a4[26][18] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][19]$_SDFFE_PP0P_  (.D(_00922_),
    .Q(\core.CPU_Xreg_value_a4[26][19] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][1]$_SDFFE_PP1P_  (.D(_00923_),
    .Q(\core.CPU_Xreg_value_a4[26][1] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][20]$_SDFFE_PP0P_  (.D(_00924_),
    .Q(\core.CPU_Xreg_value_a4[26][20] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][21]$_SDFFE_PP0P_  (.D(_00925_),
    .Q(\core.CPU_Xreg_value_a4[26][21] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][22]$_SDFFE_PP0P_  (.D(_00926_),
    .Q(\core.CPU_Xreg_value_a4[26][22] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][23]$_SDFFE_PP0P_  (.D(_00927_),
    .Q(\core.CPU_Xreg_value_a4[26][23] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][24]$_SDFFE_PP0P_  (.D(_00928_),
    .Q(\core.CPU_Xreg_value_a4[26][24] ),
    .CLK(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][25]$_SDFFE_PP0P_  (.D(_00929_),
    .Q(\core.CPU_Xreg_value_a4[26][25] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][26]$_SDFFE_PP0P_  (.D(_00930_),
    .Q(\core.CPU_Xreg_value_a4[26][26] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][27]$_SDFFE_PP0P_  (.D(_00931_),
    .Q(\core.CPU_Xreg_value_a4[26][27] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][28]$_SDFFE_PP0P_  (.D(_00932_),
    .Q(\core.CPU_Xreg_value_a4[26][28] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][29]$_SDFFE_PP0P_  (.D(_00933_),
    .Q(\core.CPU_Xreg_value_a4[26][29] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][2]$_SDFFE_PP0P_  (.D(_00934_),
    .Q(\core.CPU_Xreg_value_a4[26][2] ),
    .CLK(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][30]$_SDFFE_PP0P_  (.D(_00935_),
    .Q(\core.CPU_Xreg_value_a4[26][30] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][31]$_SDFFE_PP0P_  (.D(_00936_),
    .Q(\core.CPU_Xreg_value_a4[26][31] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][3]$_SDFFE_PP1P_  (.D(_00937_),
    .Q(\core.CPU_Xreg_value_a4[26][3] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][4]$_SDFFE_PP1P_  (.D(_00938_),
    .Q(\core.CPU_Xreg_value_a4[26][4] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][5]$_SDFFE_PP0P_  (.D(_00939_),
    .Q(\core.CPU_Xreg_value_a4[26][5] ),
    .CLK(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][6]$_SDFFE_PP0P_  (.D(_00940_),
    .Q(\core.CPU_Xreg_value_a4[26][6] ),
    .CLK(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][7]$_SDFFE_PP0P_  (.D(_00941_),
    .Q(\core.CPU_Xreg_value_a4[26][7] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][8]$_SDFFE_PP0P_  (.D(_00942_),
    .Q(\core.CPU_Xreg_value_a4[26][8] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[26][9]$_SDFFE_PP0P_  (.D(_00943_),
    .Q(\core.CPU_Xreg_value_a4[26][9] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][0]$_SDFFE_PP1P_  (.D(_00944_),
    .Q(\core.CPU_Xreg_value_a4[27][0] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][10]$_SDFFE_PP0P_  (.D(_00945_),
    .Q(\core.CPU_Xreg_value_a4[27][10] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][11]$_SDFFE_PP0P_  (.D(_00946_),
    .Q(\core.CPU_Xreg_value_a4[27][11] ),
    .CLK(clknet_leaf_110_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][12]$_SDFFE_PP0P_  (.D(_00947_),
    .Q(\core.CPU_Xreg_value_a4[27][12] ),
    .CLK(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][13]$_SDFFE_PP0P_  (.D(_00948_),
    .Q(\core.CPU_Xreg_value_a4[27][13] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][14]$_SDFFE_PP0P_  (.D(_00949_),
    .Q(\core.CPU_Xreg_value_a4[27][14] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][15]$_SDFFE_PP0P_  (.D(_00950_),
    .Q(\core.CPU_Xreg_value_a4[27][15] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][16]$_SDFFE_PP0P_  (.D(_00951_),
    .Q(\core.CPU_Xreg_value_a4[27][16] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][17]$_SDFFE_PP0P_  (.D(_00952_),
    .Q(\core.CPU_Xreg_value_a4[27][17] ),
    .CLK(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][18]$_SDFFE_PP0P_  (.D(_00953_),
    .Q(\core.CPU_Xreg_value_a4[27][18] ),
    .CLK(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][19]$_SDFFE_PP0P_  (.D(_00954_),
    .Q(\core.CPU_Xreg_value_a4[27][19] ),
    .CLK(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][1]$_SDFFE_PP1P_  (.D(_00955_),
    .Q(\core.CPU_Xreg_value_a4[27][1] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][20]$_SDFFE_PP0P_  (.D(_00956_),
    .Q(\core.CPU_Xreg_value_a4[27][20] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][21]$_SDFFE_PP0P_  (.D(_00957_),
    .Q(\core.CPU_Xreg_value_a4[27][21] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][22]$_SDFFE_PP0P_  (.D(_00958_),
    .Q(\core.CPU_Xreg_value_a4[27][22] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][23]$_SDFFE_PP0P_  (.D(_00959_),
    .Q(\core.CPU_Xreg_value_a4[27][23] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][24]$_SDFFE_PP0P_  (.D(_00960_),
    .Q(\core.CPU_Xreg_value_a4[27][24] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][25]$_SDFFE_PP0P_  (.D(_00961_),
    .Q(\core.CPU_Xreg_value_a4[27][25] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][26]$_SDFFE_PP0P_  (.D(_00962_),
    .Q(\core.CPU_Xreg_value_a4[27][26] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][27]$_SDFFE_PP0P_  (.D(_00963_),
    .Q(\core.CPU_Xreg_value_a4[27][27] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][28]$_SDFFE_PP0P_  (.D(_00964_),
    .Q(\core.CPU_Xreg_value_a4[27][28] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][29]$_SDFFE_PP0P_  (.D(_00965_),
    .Q(\core.CPU_Xreg_value_a4[27][29] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][2]$_SDFFE_PP0P_  (.D(_00966_),
    .Q(\core.CPU_Xreg_value_a4[27][2] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][30]$_SDFFE_PP0P_  (.D(_00967_),
    .Q(\core.CPU_Xreg_value_a4[27][30] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][31]$_SDFFE_PP0P_  (.D(_00968_),
    .Q(\core.CPU_Xreg_value_a4[27][31] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][3]$_SDFFE_PP1P_  (.D(_00969_),
    .Q(\core.CPU_Xreg_value_a4[27][3] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][4]$_SDFFE_PP1P_  (.D(_00970_),
    .Q(\core.CPU_Xreg_value_a4[27][4] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][5]$_SDFFE_PP0P_  (.D(_00971_),
    .Q(\core.CPU_Xreg_value_a4[27][5] ),
    .CLK(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][6]$_SDFFE_PP0P_  (.D(_00972_),
    .Q(\core.CPU_Xreg_value_a4[27][6] ),
    .CLK(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][7]$_SDFFE_PP0P_  (.D(_00973_),
    .Q(\core.CPU_Xreg_value_a4[27][7] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][8]$_SDFFE_PP0P_  (.D(_00974_),
    .Q(\core.CPU_Xreg_value_a4[27][8] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[27][9]$_SDFFE_PP0P_  (.D(_00975_),
    .Q(\core.CPU_Xreg_value_a4[27][9] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][0]$_SDFFE_PP0P_  (.D(_00976_),
    .Q(\core.CPU_Xreg_value_a4[2][0] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][10]$_SDFFE_PP0P_  (.D(_00977_),
    .Q(\core.CPU_Xreg_value_a4[2][10] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][11]$_SDFFE_PP0P_  (.D(_00978_),
    .Q(\core.CPU_Xreg_value_a4[2][11] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][12]$_SDFFE_PP0P_  (.D(_00979_),
    .Q(\core.CPU_Xreg_value_a4[2][12] ),
    .CLK(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][13]$_SDFFE_PP0P_  (.D(_00980_),
    .Q(\core.CPU_Xreg_value_a4[2][13] ),
    .CLK(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][14]$_SDFFE_PP0P_  (.D(_00981_),
    .Q(\core.CPU_Xreg_value_a4[2][14] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][15]$_SDFFE_PP0P_  (.D(_00982_),
    .Q(\core.CPU_Xreg_value_a4[2][15] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][16]$_SDFFE_PP0P_  (.D(_00983_),
    .Q(\core.CPU_Xreg_value_a4[2][16] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][17]$_SDFFE_PP0P_  (.D(_00984_),
    .Q(\core.CPU_Xreg_value_a4[2][17] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][18]$_SDFFE_PP0P_  (.D(_00985_),
    .Q(\core.CPU_Xreg_value_a4[2][18] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][19]$_SDFFE_PP0P_  (.D(_00986_),
    .Q(\core.CPU_Xreg_value_a4[2][19] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][1]$_SDFFE_PP1P_  (.D(_00987_),
    .Q(\core.CPU_Xreg_value_a4[2][1] ),
    .CLK(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][20]$_SDFFE_PP0P_  (.D(_00988_),
    .Q(\core.CPU_Xreg_value_a4[2][20] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][21]$_SDFFE_PP0P_  (.D(_00989_),
    .Q(\core.CPU_Xreg_value_a4[2][21] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][22]$_SDFFE_PP0P_  (.D(_00990_),
    .Q(\core.CPU_Xreg_value_a4[2][22] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][23]$_SDFFE_PP0P_  (.D(_00991_),
    .Q(\core.CPU_Xreg_value_a4[2][23] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][24]$_SDFFE_PP0P_  (.D(_00992_),
    .Q(\core.CPU_Xreg_value_a4[2][24] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][25]$_SDFFE_PP0P_  (.D(_00993_),
    .Q(\core.CPU_Xreg_value_a4[2][25] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][26]$_SDFFE_PP0P_  (.D(_00994_),
    .Q(\core.CPU_Xreg_value_a4[2][26] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][27]$_SDFFE_PP0P_  (.D(_00995_),
    .Q(\core.CPU_Xreg_value_a4[2][27] ),
    .CLK(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][28]$_SDFFE_PP0P_  (.D(_00996_),
    .Q(\core.CPU_Xreg_value_a4[2][28] ),
    .CLK(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][29]$_SDFFE_PP0P_  (.D(_00997_),
    .Q(\core.CPU_Xreg_value_a4[2][29] ),
    .CLK(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][2]$_SDFFE_PP0P_  (.D(_00998_),
    .Q(\core.CPU_Xreg_value_a4[2][2] ),
    .CLK(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][30]$_SDFFE_PP0P_  (.D(_00999_),
    .Q(\core.CPU_Xreg_value_a4[2][30] ),
    .CLK(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][31]$_SDFFE_PP0P_  (.D(_01000_),
    .Q(\core.CPU_Xreg_value_a4[2][31] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][3]$_SDFFE_PP0P_  (.D(_01001_),
    .Q(\core.CPU_Xreg_value_a4[2][3] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][4]$_SDFFE_PP0P_  (.D(_01002_),
    .Q(\core.CPU_Xreg_value_a4[2][4] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][5]$_SDFFE_PP0P_  (.D(_01003_),
    .Q(\core.CPU_Xreg_value_a4[2][5] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][6]$_SDFFE_PP0P_  (.D(_01004_),
    .Q(\core.CPU_Xreg_value_a4[2][6] ),
    .CLK(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][7]$_SDFFE_PP0P_  (.D(_01005_),
    .Q(\core.CPU_Xreg_value_a4[2][7] ),
    .CLK(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][8]$_SDFFE_PP0P_  (.D(_01006_),
    .Q(\core.CPU_Xreg_value_a4[2][8] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[2][9]$_SDFFE_PP0P_  (.D(_01007_),
    .Q(\core.CPU_Xreg_value_a4[2][9] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][0]$_SDFFE_PP1P_  (.D(_01008_),
    .Q(\core.CPU_Xreg_value_a4[3][0] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][10]$_SDFFE_PP0P_  (.D(_01009_),
    .Q(\core.CPU_Xreg_value_a4[3][10] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][11]$_SDFFE_PP0P_  (.D(_01010_),
    .Q(\core.CPU_Xreg_value_a4[3][11] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][12]$_SDFFE_PP0P_  (.D(_01011_),
    .Q(\core.CPU_Xreg_value_a4[3][12] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][13]$_SDFFE_PP0P_  (.D(_01012_),
    .Q(\core.CPU_Xreg_value_a4[3][13] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][14]$_SDFFE_PP0P_  (.D(_01013_),
    .Q(\core.CPU_Xreg_value_a4[3][14] ),
    .CLK(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][15]$_SDFFE_PP0P_  (.D(_01014_),
    .Q(\core.CPU_Xreg_value_a4[3][15] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][16]$_SDFFE_PP0P_  (.D(_01015_),
    .Q(\core.CPU_Xreg_value_a4[3][16] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][17]$_SDFFE_PP0P_  (.D(_01016_),
    .Q(\core.CPU_Xreg_value_a4[3][17] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][18]$_SDFFE_PP0P_  (.D(_01017_),
    .Q(\core.CPU_Xreg_value_a4[3][18] ),
    .CLK(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][19]$_SDFFE_PP0P_  (.D(_01018_),
    .Q(\core.CPU_Xreg_value_a4[3][19] ),
    .CLK(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][1]$_SDFFE_PP1P_  (.D(_01019_),
    .Q(\core.CPU_Xreg_value_a4[3][1] ),
    .CLK(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][20]$_SDFFE_PP0P_  (.D(_01020_),
    .Q(\core.CPU_Xreg_value_a4[3][20] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][21]$_SDFFE_PP0P_  (.D(_01021_),
    .Q(\core.CPU_Xreg_value_a4[3][21] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][22]$_SDFFE_PP0P_  (.D(_01022_),
    .Q(\core.CPU_Xreg_value_a4[3][22] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][23]$_SDFFE_PP0P_  (.D(_01023_),
    .Q(\core.CPU_Xreg_value_a4[3][23] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][24]$_SDFFE_PP0P_  (.D(_01024_),
    .Q(\core.CPU_Xreg_value_a4[3][24] ),
    .CLK(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][25]$_SDFFE_PP0P_  (.D(_01025_),
    .Q(\core.CPU_Xreg_value_a4[3][25] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][26]$_SDFFE_PP0P_  (.D(_01026_),
    .Q(\core.CPU_Xreg_value_a4[3][26] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][27]$_SDFFE_PP0P_  (.D(_01027_),
    .Q(\core.CPU_Xreg_value_a4[3][27] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][28]$_SDFFE_PP0P_  (.D(_01028_),
    .Q(\core.CPU_Xreg_value_a4[3][28] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][29]$_SDFFE_PP0P_  (.D(_01029_),
    .Q(\core.CPU_Xreg_value_a4[3][29] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][2]$_SDFFE_PP0P_  (.D(_01030_),
    .Q(\core.CPU_Xreg_value_a4[3][2] ),
    .CLK(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][30]$_SDFFE_PP0P_  (.D(_01031_),
    .Q(\core.CPU_Xreg_value_a4[3][30] ),
    .CLK(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][31]$_SDFFE_PP0P_  (.D(_01032_),
    .Q(\core.CPU_Xreg_value_a4[3][31] ),
    .CLK(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][3]$_SDFFE_PP0P_  (.D(_01033_),
    .Q(\core.CPU_Xreg_value_a4[3][3] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][4]$_SDFFE_PP0P_  (.D(_01034_),
    .Q(\core.CPU_Xreg_value_a4[3][4] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][5]$_SDFFE_PP0P_  (.D(_01035_),
    .Q(\core.CPU_Xreg_value_a4[3][5] ),
    .CLK(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][6]$_SDFFE_PP0P_  (.D(_01036_),
    .Q(\core.CPU_Xreg_value_a4[3][6] ),
    .CLK(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][7]$_SDFFE_PP0P_  (.D(_01037_),
    .Q(\core.CPU_Xreg_value_a4[3][7] ),
    .CLK(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][8]$_SDFFE_PP0P_  (.D(_01038_),
    .Q(\core.CPU_Xreg_value_a4[3][8] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[3][9]$_SDFFE_PP0P_  (.D(_01039_),
    .Q(\core.CPU_Xreg_value_a4[3][9] ),
    .CLK(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][0]$_SDFFE_PP0P_  (.D(_01040_),
    .Q(\core.CPU_Xreg_value_a4[8][0] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][10]$_SDFFE_PP0P_  (.D(_01041_),
    .Q(\core.CPU_Xreg_value_a4[8][10] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][11]$_SDFFE_PP0P_  (.D(_01042_),
    .Q(\core.CPU_Xreg_value_a4[8][11] ),
    .CLK(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][12]$_SDFFE_PP0P_  (.D(_01043_),
    .Q(\core.CPU_Xreg_value_a4[8][12] ),
    .CLK(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][13]$_SDFFE_PP0P_  (.D(_01044_),
    .Q(\core.CPU_Xreg_value_a4[8][13] ),
    .CLK(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][14]$_SDFFE_PP0P_  (.D(_01045_),
    .Q(\core.CPU_Xreg_value_a4[8][14] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][15]$_SDFFE_PP0P_  (.D(_01046_),
    .Q(\core.CPU_Xreg_value_a4[8][15] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][16]$_SDFFE_PP0P_  (.D(_01047_),
    .Q(\core.CPU_Xreg_value_a4[8][16] ),
    .CLK(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][17]$_SDFFE_PP0P_  (.D(_01048_),
    .Q(\core.CPU_Xreg_value_a4[8][17] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][18]$_SDFFE_PP0P_  (.D(_01049_),
    .Q(\core.CPU_Xreg_value_a4[8][18] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][19]$_SDFFE_PP0P_  (.D(_01050_),
    .Q(\core.CPU_Xreg_value_a4[8][19] ),
    .CLK(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][1]$_SDFFE_PP0P_  (.D(_01051_),
    .Q(\core.CPU_Xreg_value_a4[8][1] ),
    .CLK(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][20]$_SDFFE_PP0P_  (.D(_01052_),
    .Q(\core.CPU_Xreg_value_a4[8][20] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][21]$_SDFFE_PP0P_  (.D(_01053_),
    .Q(\core.CPU_Xreg_value_a4[8][21] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][22]$_SDFFE_PP0P_  (.D(_01054_),
    .Q(\core.CPU_Xreg_value_a4[8][22] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][23]$_SDFFE_PP0P_  (.D(_01055_),
    .Q(\core.CPU_Xreg_value_a4[8][23] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][24]$_SDFFE_PP0P_  (.D(_01056_),
    .Q(\core.CPU_Xreg_value_a4[8][24] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][25]$_SDFFE_PP0P_  (.D(_01057_),
    .Q(\core.CPU_Xreg_value_a4[8][25] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][26]$_SDFFE_PP0P_  (.D(_01058_),
    .Q(\core.CPU_Xreg_value_a4[8][26] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][27]$_SDFFE_PP0P_  (.D(_01059_),
    .Q(\core.CPU_Xreg_value_a4[8][27] ),
    .CLK(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][28]$_SDFFE_PP0P_  (.D(_01060_),
    .Q(\core.CPU_Xreg_value_a4[8][28] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][29]$_SDFFE_PP0P_  (.D(_01061_),
    .Q(\core.CPU_Xreg_value_a4[8][29] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][2]$_SDFFE_PP0P_  (.D(_01062_),
    .Q(\core.CPU_Xreg_value_a4[8][2] ),
    .CLK(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][30]$_SDFFE_PP0P_  (.D(_01063_),
    .Q(\core.CPU_Xreg_value_a4[8][30] ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][31]$_SDFFE_PP0P_  (.D(_01064_),
    .Q(\core.CPU_Xreg_value_a4[8][31] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][3]$_SDFFE_PP1P_  (.D(_01065_),
    .Q(\core.CPU_Xreg_value_a4[8][3] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][4]$_SDFFE_PP0P_  (.D(_01066_),
    .Q(\core.CPU_Xreg_value_a4[8][4] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][5]$_SDFFE_PP0P_  (.D(_01067_),
    .Q(\core.CPU_Xreg_value_a4[8][5] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][6]$_SDFFE_PP0P_  (.D(_01068_),
    .Q(\core.CPU_Xreg_value_a4[8][6] ),
    .CLK(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][7]$_SDFFE_PP0P_  (.D(_01069_),
    .Q(\core.CPU_Xreg_value_a4[8][7] ),
    .CLK(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][8]$_SDFFE_PP0P_  (.D(_01070_),
    .Q(\core.CPU_Xreg_value_a4[8][8] ),
    .CLK(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[8][9]$_SDFFE_PP0P_  (.D(_01071_),
    .Q(\core.CPU_Xreg_value_a4[8][9] ),
    .CLK(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][0]$_SDFFE_PP1P_  (.D(_01072_),
    .Q(\core.CPU_Xreg_value_a4[9][0] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][10]$_SDFFE_PP0P_  (.D(_01073_),
    .Q(\core.CPU_Xreg_value_a4[9][10] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][11]$_SDFFE_PP0P_  (.D(_01074_),
    .Q(\core.CPU_Xreg_value_a4[9][11] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][12]$_SDFFE_PP0P_  (.D(_01075_),
    .Q(\core.CPU_Xreg_value_a4[9][12] ),
    .CLK(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][13]$_SDFFE_PP0P_  (.D(_01076_),
    .Q(\core.CPU_Xreg_value_a4[9][13] ),
    .CLK(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][14]$_SDFFE_PP0P_  (.D(_01077_),
    .Q(\core.CPU_Xreg_value_a4[9][14] ),
    .CLK(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][15]$_SDFFE_PP0P_  (.D(_01078_),
    .Q(\core.CPU_Xreg_value_a4[9][15] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][16]$_SDFFE_PP0P_  (.D(_01079_),
    .Q(\core.CPU_Xreg_value_a4[9][16] ),
    .CLK(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][17]$_SDFFE_PP0P_  (.D(_01080_),
    .Q(\core.CPU_Xreg_value_a4[9][17] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][18]$_SDFFE_PP0P_  (.D(_01081_),
    .Q(\core.CPU_Xreg_value_a4[9][18] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][19]$_SDFFE_PP0P_  (.D(_01082_),
    .Q(\core.CPU_Xreg_value_a4[9][19] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][1]$_SDFFE_PP0P_  (.D(_01083_),
    .Q(\core.CPU_Xreg_value_a4[9][1] ),
    .CLK(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][20]$_SDFFE_PP0P_  (.D(_01084_),
    .Q(\core.CPU_Xreg_value_a4[9][20] ),
    .CLK(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][21]$_SDFFE_PP0P_  (.D(_01085_),
    .Q(\core.CPU_Xreg_value_a4[9][21] ),
    .CLK(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][22]$_SDFFE_PP0P_  (.D(_01086_),
    .Q(\core.CPU_Xreg_value_a4[9][22] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][23]$_SDFFE_PP0P_  (.D(_01087_),
    .Q(\core.CPU_Xreg_value_a4[9][23] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][24]$_SDFFE_PP0P_  (.D(_01088_),
    .Q(\core.CPU_Xreg_value_a4[9][24] ),
    .CLK(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][25]$_SDFFE_PP0P_  (.D(_01089_),
    .Q(\core.CPU_Xreg_value_a4[9][25] ),
    .CLK(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][26]$_SDFFE_PP0P_  (.D(_01090_),
    .Q(\core.CPU_Xreg_value_a4[9][26] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][27]$_SDFFE_PP0P_  (.D(_01091_),
    .Q(\core.CPU_Xreg_value_a4[9][27] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][28]$_SDFFE_PP0P_  (.D(_01092_),
    .Q(\core.CPU_Xreg_value_a4[9][28] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][29]$_SDFFE_PP0P_  (.D(_01093_),
    .Q(\core.CPU_Xreg_value_a4[9][29] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][2]$_SDFFE_PP0P_  (.D(_01094_),
    .Q(\core.CPU_Xreg_value_a4[9][2] ),
    .CLK(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][30]$_SDFFE_PP0P_  (.D(_01095_),
    .Q(\core.CPU_Xreg_value_a4[9][30] ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][31]$_SDFFE_PP0P_  (.D(_01096_),
    .Q(\core.CPU_Xreg_value_a4[9][31] ),
    .CLK(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][3]$_SDFFE_PP1P_  (.D(_01097_),
    .Q(\core.CPU_Xreg_value_a4[9][3] ),
    .CLK(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][4]$_SDFFE_PP0P_  (.D(_01098_),
    .Q(\core.CPU_Xreg_value_a4[9][4] ),
    .CLK(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][5]$_SDFFE_PP0P_  (.D(_01099_),
    .Q(\core.CPU_Xreg_value_a4[9][5] ),
    .CLK(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][6]$_SDFFE_PP0P_  (.D(_01100_),
    .Q(\core.CPU_Xreg_value_a4[9][6] ),
    .CLK(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][7]$_SDFFE_PP0P_  (.D(_01101_),
    .Q(\core.CPU_Xreg_value_a4[9][7] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][8]$_SDFFE_PP0P_  (.D(_01102_),
    .Q(\core.CPU_Xreg_value_a4[9][8] ),
    .CLK(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a4[9][9]$_SDFFE_PP0P_  (.D(_01103_),
    .Q(\core.CPU_Xreg_value_a4[9][9] ),
    .CLK(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][0]$_DFF_P_  (.D(net620),
    .Q(\core.CPU_Xreg_value_a5[17][0] ),
    .CLK(clknet_leaf_112_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][1]$_DFF_P_  (.D(net619),
    .Q(\core.CPU_Xreg_value_a5[17][1] ),
    .CLK(clknet_leaf_112_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][2]$_DFF_P_  (.D(net618),
    .Q(\core.CPU_Xreg_value_a5[17][2] ),
    .CLK(clknet_leaf_111_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][3]$_DFF_P_  (.D(\core.CPU_Xreg_value_a4[17][3] ),
    .Q(\core.CPU_Xreg_value_a5[17][3] ),
    .CLK(clknet_leaf_111_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][4]$_DFF_P_  (.D(net617),
    .Q(\core.CPU_Xreg_value_a5[17][4] ),
    .CLK(clknet_leaf_111_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][5]$_DFF_P_  (.D(net616),
    .Q(\core.CPU_Xreg_value_a5[17][5] ),
    .CLK(clknet_leaf_111_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][6]$_DFF_P_  (.D(\core.CPU_Xreg_value_a4[17][6] ),
    .Q(\core.CPU_Xreg_value_a5[17][6] ),
    .CLK(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][7]$_DFF_P_  (.D(\core.CPU_Xreg_value_a4[17][7] ),
    .Q(\core.CPU_Xreg_value_a5[17][7] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][8]$_DFF_P_  (.D(\core.CPU_Xreg_value_a4[17][8] ),
    .Q(\core.CPU_Xreg_value_a5[17][8] ),
    .CLK(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_Xreg_value_a5[17][9]$_DFF_P_  (.D(\core.CPU_Xreg_value_a4[17][9] ),
    .Q(\core.CPU_Xreg_value_a5[17][9] ),
    .CLK(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_br_tgt_pc_a3[0]$_DFF_P_  (.D(\core.CPU_br_tgt_pc_a2[0] ),
    .Q(\core.CPU_br_tgt_pc_a3[0] ),
    .CLK(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_br_tgt_pc_a3[1]$_DFF_P_  (.D(\core.CPU_br_tgt_pc_a2[1] ),
    .Q(\core.CPU_br_tgt_pc_a3[1] ),
    .CLK(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_br_tgt_pc_a3[2]$_DFF_P_  (.D(\core.CPU_br_tgt_pc_a2[2] ),
    .Q(\core.CPU_br_tgt_pc_a3[2] ),
    .CLK(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_br_tgt_pc_a3[3]$_DFF_P_  (.D(\core.CPU_br_tgt_pc_a2[3] ),
    .Q(\core.CPU_br_tgt_pc_a3[3] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_br_tgt_pc_a3[4]$_DFF_P_  (.D(\core.CPU_br_tgt_pc_a2[4] ),
    .Q(\core.CPU_br_tgt_pc_a3[4] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_br_tgt_pc_a3[5]$_DFF_P_  (.D(\core.CPU_br_tgt_pc_a2[5] ),
    .Q(\core.CPU_br_tgt_pc_a3[5] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[0]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[0] ),
    .Q(\core.CPU_dmem_rd_data_a5[0] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[10]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[10] ),
    .Q(\core.CPU_dmem_rd_data_a5[10] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[11]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[11] ),
    .Q(\core.CPU_dmem_rd_data_a5[11] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[12]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[12] ),
    .Q(\core.CPU_dmem_rd_data_a5[12] ),
    .CLK(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[13]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[13] ),
    .Q(\core.CPU_dmem_rd_data_a5[13] ),
    .CLK(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[14]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[14] ),
    .Q(\core.CPU_dmem_rd_data_a5[14] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[15]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[15] ),
    .Q(\core.CPU_dmem_rd_data_a5[15] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[16]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[16] ),
    .Q(\core.CPU_dmem_rd_data_a5[16] ),
    .CLK(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[17]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[17] ),
    .Q(\core.CPU_dmem_rd_data_a5[17] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[18]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[18] ),
    .Q(\core.CPU_dmem_rd_data_a5[18] ),
    .CLK(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[19]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[19] ),
    .Q(\core.CPU_dmem_rd_data_a5[19] ),
    .CLK(clknet_leaf_68_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[1]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[1] ),
    .Q(\core.CPU_dmem_rd_data_a5[1] ),
    .CLK(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[20]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[20] ),
    .Q(\core.CPU_dmem_rd_data_a5[20] ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[21]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[21] ),
    .Q(\core.CPU_dmem_rd_data_a5[21] ),
    .CLK(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[22]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[22] ),
    .Q(\core.CPU_dmem_rd_data_a5[22] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[23]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[23] ),
    .Q(\core.CPU_dmem_rd_data_a5[23] ),
    .CLK(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[24]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[24] ),
    .Q(\core.CPU_dmem_rd_data_a5[24] ),
    .CLK(clknet_leaf_66_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[25]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[25] ),
    .Q(\core.CPU_dmem_rd_data_a5[25] ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[26]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[26] ),
    .Q(\core.CPU_dmem_rd_data_a5[26] ),
    .CLK(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[27]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[27] ),
    .Q(\core.CPU_dmem_rd_data_a5[27] ),
    .CLK(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[28]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[28] ),
    .Q(\core.CPU_dmem_rd_data_a5[28] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[29]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[29] ),
    .Q(\core.CPU_dmem_rd_data_a5[29] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[2]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[2] ),
    .Q(\core.CPU_dmem_rd_data_a5[2] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[30]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[30] ),
    .Q(\core.CPU_dmem_rd_data_a5[30] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[31]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[31] ),
    .Q(\core.CPU_dmem_rd_data_a5[31] ),
    .CLK(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[3]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[3] ),
    .Q(\core.CPU_dmem_rd_data_a5[3] ),
    .CLK(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[4]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[4] ),
    .Q(\core.CPU_dmem_rd_data_a5[4] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[5]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[5] ),
    .Q(\core.CPU_dmem_rd_data_a5[5] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[6]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[6] ),
    .Q(\core.CPU_dmem_rd_data_a5[6] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[7]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[7] ),
    .Q(\core.CPU_dmem_rd_data_a5[7] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[8]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[8] ),
    .Q(\core.CPU_dmem_rd_data_a5[8] ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_dmem_rd_data_a5[9]$_DFF_P_  (.D(\core.w_CPU_dmem_rd_data_a4[9] ),
    .Q(\core.CPU_dmem_rd_data_a5[9] ),
    .CLK(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imem_rd_addr_a1[0]$_SDFF_PP0_  (.D(_01104_),
    .Q(\core.CPU_imem_rd_addr_a1[0] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imem_rd_addr_a1[1]$_SDFF_PP0_  (.D(_01105_),
    .Q(\core.CPU_imem_rd_addr_a1[1] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imem_rd_addr_a1[2]$_SDFF_PP0_  (.D(_01106_),
    .Q(\core.CPU_imem_rd_addr_a1[2] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imem_rd_addr_a1[3]$_SDFF_PP0_  (.D(_01107_),
    .Q(\core.CPU_imem_rd_addr_a1[3] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a2[0]$_DFF_P_  (.D(\core.CPU_imm_a1[0] ),
    .Q(\core.CPU_imm_a2[0] ),
    .CLK(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a2[10]$_DFF_P_  (.D(\core.CPU_imm_a1[10] ),
    .Q(\core.CPU_imm_a2[10] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a2[11]$_DFF_P_  (.D(\core.CPU_imm_a1[11] ),
    .Q(\core.CPU_imm_a2[11] ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a2[1]$_DFF_P_  (.D(\core.CPU_imm_a1[1] ),
    .Q(\core.CPU_imm_a2[1] ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a2[30]$_DFF_P_  (.D(\core.CPU_imm_a1[12] ),
    .Q(\core.CPU_imm_a2[12] ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a2[3]$_DFF_P_  (.D(\core.CPU_imm_a1[3] ),
    .Q(\core.CPU_imm_a2[3] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a2[4]$_SDFF_PP0_  (.D(_01108_),
    .Q(\core.CPU_imm_a2[4] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a2[5]$_DFF_P_  (.D(\core.CPU_imm_a1[5] ),
    .Q(\core.CPU_imm_a2[5] ),
    .CLK(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a3[0]$_DFF_P_  (.D(\core.CPU_imm_a2[0] ),
    .Q(\core.CPU_imm_a3[0] ),
    .CLK(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a3[10]$_DFF_P_  (.D(\core.CPU_imm_a2[10] ),
    .Q(\core.CPU_imm_a3[10] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a3[11]$_DFF_P_  (.D(\core.CPU_imm_a2[11] ),
    .Q(\core.CPU_imm_a3[11] ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a3[1]$_DFF_P_  (.D(\core.CPU_imm_a2[1] ),
    .Q(\core.CPU_imm_a3[1] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a3[30]$_DFF_P_  (.D(\core.CPU_imm_a2[12] ),
    .Q(\core.CPU_imm_a3[12] ),
    .CLK(clknet_leaf_68_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a3[3]$_DFF_P_  (.D(\core.CPU_imm_a2[3] ),
    .Q(\core.CPU_imm_a3[3] ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a3[4]$_DFF_P_  (.D(\core.CPU_imm_a2[4] ),
    .Q(\core.CPU_imm_a3[4] ),
    .CLK(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_imm_a3[5]$_DFF_P_  (.D(\core.CPU_imm_a2[5] ),
    .Q(\core.CPU_imm_a3[5] ),
    .CLK(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a2[0]$_DFF_P_  (.D(\core.CPU_inc_pc_a1[0] ),
    .Q(\core.CPU_inc_pc_a2[0] ),
    .CLK(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a2[1]$_DFF_P_  (.D(\core.CPU_inc_pc_a1[1] ),
    .Q(\core.CPU_inc_pc_a2[1] ),
    .CLK(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a2[2]$_DFF_P_  (.D(\core.CPU_inc_pc_a1[2] ),
    .Q(\core.CPU_inc_pc_a2[2] ),
    .CLK(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a2[3]$_DFF_P_  (.D(\core.CPU_inc_pc_a1[3] ),
    .Q(\core.CPU_inc_pc_a2[3] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a2[4]$_DFF_P_  (.D(\core.CPU_inc_pc_a1[4] ),
    .Q(\core.CPU_inc_pc_a2[4] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a2[5]$_DFF_P_  (.D(\core.CPU_inc_pc_a1[5] ),
    .Q(\core.CPU_inc_pc_a2[5] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a3[0]$_DFF_P_  (.D(\core.CPU_inc_pc_a2[0] ),
    .Q(\core.CPU_inc_pc_a3[0] ),
    .CLK(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a3[1]$_DFF_P_  (.D(\core.CPU_inc_pc_a2[1] ),
    .Q(\core.CPU_inc_pc_a3[1] ),
    .CLK(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a3[2]$_DFF_P_  (.D(\core.CPU_inc_pc_a2[2] ),
    .Q(\core.CPU_inc_pc_a3[2] ),
    .CLK(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a3[3]$_DFF_P_  (.D(\core.CPU_inc_pc_a2[3] ),
    .Q(\core.CPU_inc_pc_a3[3] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a3[4]$_DFF_P_  (.D(\core.CPU_inc_pc_a2[4] ),
    .Q(\core.CPU_inc_pc_a3[4] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_inc_pc_a3[5]$_DFF_P_  (.D(\core.CPU_inc_pc_a2[5] ),
    .Q(\core.CPU_inc_pc_a3[5] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_add_a2$_DFF_P_  (.D(\core.CPU_is_add_a1 ),
    .Q(\core.CPU_is_add_a2 ),
    .CLK(clknet_leaf_68_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_add_a3$_DFF_P_  (.D(\core.CPU_is_add_a2 ),
    .Q(\core.CPU_is_add_a3 ),
    .CLK(clknet_leaf_68_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_addi_a2$_DFF_P_  (.D(\core.CPU_is_addi_a1 ),
    .Q(\core.CPU_is_addi_a2 ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_2 \core.CPU_is_addi_a3$_DFF_P_  (.D(\core.CPU_is_addi_a2 ),
    .Q(\core.CPU_is_addi_a3 ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_beq_a2$_DFF_P_  (.D(\core.CPU_is_beq_a1 ),
    .Q(\core.CPU_is_beq_a2 ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_beq_a3$_DFF_P_  (.D(\core.CPU_is_beq_a2 ),
    .Q(\core.CPU_is_beq_a3 ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_bne_a2$_DFF_P_  (.D(\core.CPU_is_bne_a1 ),
    .Q(\core.CPU_is_bne_a2 ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_bne_a3$_DFF_P_  (.D(\core.CPU_is_bne_a2 ),
    .Q(\core.CPU_is_bne_a3 ),
    .CLK(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_load_a2$_DFF_P_  (.D(net),
    .Q(\core.CPU_is_load_a2 ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_load_a3$_DFF_P_  (.D(\core.CPU_is_load_a2 ),
    .Q(\core.CPU_is_load_a3 ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_s_instr_a2$_DFF_P_  (.D(net1),
    .Q(\core.CPU_is_s_instr_a2 ),
    .CLK(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_s_instr_a3$_DFF_P_  (.D(\core.CPU_is_s_instr_a2 ),
    .Q(\core.CPU_is_s_instr_a3 ),
    .CLK(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_s_instr_a4$_DFF_P_  (.D(\core.CPU_is_s_instr_a3 ),
    .Q(\core.CPU_is_s_instr_a4 ),
    .CLK(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_sll_a2$_DFF_P_  (.D(net2),
    .Q(\core.CPU_is_sll_a2 ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_sll_a3$_DFF_P_  (.D(\core.CPU_is_sll_a2 ),
    .Q(\core.CPU_is_sll_a3 ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_slli_a2$_DFF_P_  (.D(net3),
    .Q(\core.CPU_is_slli_a2 ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_slli_a3$_DFF_P_  (.D(\core.CPU_is_slli_a2 ),
    .Q(\core.CPU_is_slli_a3 ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_sub_a2$_DFF_P_  (.D(\core.CPU_is_sub_a1 ),
    .Q(\core.CPU_is_sub_a2 ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_is_sub_a3$_DFF_P_  (.D(\core.CPU_is_sub_a2 ),
    .Q(\core.CPU_is_sub_a3 ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_pc_a1[0]$_SDFFE_PP0P_  (.D(_01109_),
    .Q(\core.CPU_inc_pc_a1[0] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_pc_a1[1]$_SDFFE_PP0P_  (.D(_01110_),
    .Q(\core.CPU_inc_pc_a1[1] ),
    .CLK(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_pc_a2[2]$_DFF_P_  (.D(\core.CPU_imem_rd_addr_a1[0] ),
    .Q(\core.CPU_pc_a2[2] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_pc_a2[3]$_DFF_P_  (.D(\core.CPU_imem_rd_addr_a1[1] ),
    .Q(\core.CPU_pc_a2[3] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_pc_a2[4]$_DFF_P_  (.D(\core.CPU_imem_rd_addr_a1[2] ),
    .Q(\core.CPU_pc_a2[4] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_pc_a2[5]$_DFF_P_  (.D(net614),
    .Q(\core.CPU_pc_a2[5] ),
    .CLK(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a2[0]$_DFF_P_  (.D(\core.CPU_imem_rd_data_a1[7] ),
    .Q(\core.CPU_rd_a2[0] ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a2[1]$_DFF_P_  (.D(\core.CPU_imem_rd_data_a1[8] ),
    .Q(\core.CPU_rd_a2[1] ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a2[3]$_DFF_P_  (.D(\core.CPU_imem_rd_data_a1[10] ),
    .Q(\core.CPU_rd_a2[3] ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a2[4]$_DFF_P_  (.D(\core.CPU_imem_rd_data_a1[11] ),
    .Q(\core.CPU_rd_a2[4] ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a3[0]$_DFF_P_  (.D(\core.CPU_rd_a2[0] ),
    .Q(\core.CPU_rd_a3[0] ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a3[1]$_DFF_P_  (.D(\core.CPU_rd_a2[1] ),
    .Q(\core.CPU_rd_a3[1] ),
    .CLK(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a3[3]$_DFF_P_  (.D(\core.CPU_rd_a2[3] ),
    .Q(\core.CPU_rd_a3[3] ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a3[4]$_DFF_P_  (.D(\core.CPU_rd_a2[4] ),
    .Q(\core.CPU_rd_a3[4] ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a4[0]$_DFF_P_  (.D(\core.CPU_rd_a3[0] ),
    .Q(\core.CPU_rd_a4[0] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a4[1]$_DFF_P_  (.D(\core.CPU_rd_a3[1] ),
    .Q(\core.CPU_rd_a4[1] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a4[3]$_DFF_P_  (.D(\core.CPU_rd_a3[3] ),
    .Q(\core.CPU_rd_a4[3] ),
    .CLK(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a4[4]$_DFF_P_  (.D(\core.CPU_rd_a3[4] ),
    .Q(\core.CPU_rd_a4[4] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a5[0]$_DFF_P_  (.D(\core.CPU_rd_a4[0] ),
    .Q(\core.CPU_rd_a5[0] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a5[1]$_DFF_P_  (.D(\core.CPU_rd_a4[1] ),
    .Q(\core.CPU_rd_a5[1] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a5[3]$_DFF_P_  (.D(\core.CPU_rd_a4[3] ),
    .Q(\core.CPU_rd_a5[3] ),
    .CLK(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_a5[4]$_DFF_P_  (.D(\core.CPU_rd_a4[4] ),
    .Q(\core.CPU_rd_a5[4] ),
    .CLK(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_valid_a2$_DFF_P_  (.D(\core.CPU_rd_valid_a1 ),
    .Q(\core.CPU_rd_valid_a2 ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_rd_valid_a3$_DFF_P_  (.D(\core.CPU_rd_valid_a2 ),
    .Q(\core.CPU_rd_valid_a3 ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_reset_a1$_DFF_P_  (.D(net9),
    .Q(\core.CPU_reset_a1 ),
    .CLK(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_reset_a2$_DFF_P_  (.D(net608),
    .Q(\core.CPU_reset_a2 ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_4 \core.CPU_reset_a3$_DFF_P_  (.D(\core.CPU_reset_a2 ),
    .Q(\core.CPU_reset_a3 ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_4 \core.CPU_reset_a4$_DFF_P_  (.D(\core.CPU_reset_a3 ),
    .Q(\core.CPU_reset_a4 ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_result_a4[2]$_DFF_P_  (.D(\core.CPU_result_a3[2] ),
    .Q(\core.CPU_dmem_addr_a4[0] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_result_a4[3]$_DFF_P_  (.D(net372),
    .Q(\core.CPU_dmem_addr_a4[1] ),
    .CLK(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_result_a4[4]$_DFF_P_  (.D(\core.CPU_result_a3[4] ),
    .Q(\core.CPU_dmem_addr_a4[2] ),
    .CLK(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_result_a4[5]$_DFF_P_  (.D(\core.CPU_result_a3[5] ),
    .Q(\core.CPU_dmem_addr_a4[3] ),
    .CLK(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__dfxtp_4 \core.CPU_rs1_a2[0]$_SDFF_PP0_  (.D(_01111_),
    .Q(\core.CPU_rf_rd_index1_a2[0] ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_2 \core.CPU_rs1_a2[1]$_SDFF_PP0_  (.D(_01112_),
    .Q(\core.CPU_rf_rd_index1_a2[1] ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_4 \core.CPU_rs1_a2[4]$_SDFF_PP0_  (.D(_01113_),
    .Q(\core.CPU_rf_rd_index1_a2[4] ),
    .CLK(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__dfxtp_4 \core.CPU_rs2_a2[0]$_DFF_P_  (.D(\core.CPU_imem_rd_data_a1[20] ),
    .Q(\core.CPU_rf_rd_index2_a2[0] ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_4 \core.CPU_rs2_a2[1]$_DFF_P_  (.D(\core.CPU_imem_rd_data_a1[21] ),
    .Q(\core.CPU_rf_rd_index2_a2[1] ),
    .CLK(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__dfxtp_4 \core.CPU_rs2_a2[3]$_DFF_P_  (.D(\core.CPU_imem_rd_data_a1[23] ),
    .Q(\core.CPU_rf_rd_index2_a2[3] ),
    .CLK(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[0]$_DFF_P_  (.D(net374),
    .Q(\core.CPU_src1_value_a3[0] ),
    .CLK(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[10]$_DFF_P_  (.D(\core.CPU_src1_value_a2[10] ),
    .Q(\core.CPU_src1_value_a3[10] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[11]$_DFF_P_  (.D(\core.CPU_src1_value_a2[11] ),
    .Q(\core.CPU_src1_value_a3[11] ),
    .CLK(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[12]$_DFF_P_  (.D(\core.CPU_src1_value_a2[12] ),
    .Q(\core.CPU_src1_value_a3[12] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[13]$_DFF_P_  (.D(\core.CPU_src1_value_a2[13] ),
    .Q(\core.CPU_src1_value_a3[13] ),
    .CLK(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[14]$_DFF_P_  (.D(\core.CPU_src1_value_a2[14] ),
    .Q(\core.CPU_src1_value_a3[14] ),
    .CLK(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[15]$_DFF_P_  (.D(\core.CPU_src1_value_a2[15] ),
    .Q(\core.CPU_src1_value_a3[15] ),
    .CLK(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[16]$_DFF_P_  (.D(\core.CPU_src1_value_a2[16] ),
    .Q(\core.CPU_src1_value_a3[16] ),
    .CLK(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[17]$_DFF_P_  (.D(\core.CPU_src1_value_a2[17] ),
    .Q(\core.CPU_src1_value_a3[17] ),
    .CLK(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[18]$_DFF_P_  (.D(\core.CPU_src1_value_a2[18] ),
    .Q(\core.CPU_src1_value_a3[18] ),
    .CLK(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[19]$_DFF_P_  (.D(\core.CPU_src1_value_a2[19] ),
    .Q(\core.CPU_src1_value_a3[19] ),
    .CLK(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[1]$_DFF_P_  (.D(\core.CPU_src1_value_a2[1] ),
    .Q(\core.CPU_src1_value_a3[1] ),
    .CLK(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[20]$_DFF_P_  (.D(\core.CPU_src1_value_a2[20] ),
    .Q(\core.CPU_src1_value_a3[20] ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[21]$_DFF_P_  (.D(\core.CPU_src1_value_a2[21] ),
    .Q(\core.CPU_src1_value_a3[21] ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[22]$_DFF_P_  (.D(\core.CPU_src1_value_a2[22] ),
    .Q(\core.CPU_src1_value_a3[22] ),
    .CLK(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[23]$_DFF_P_  (.D(\core.CPU_src1_value_a2[23] ),
    .Q(\core.CPU_src1_value_a3[23] ),
    .CLK(clknet_leaf_66_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[24]$_DFF_P_  (.D(\core.CPU_src1_value_a2[24] ),
    .Q(\core.CPU_src1_value_a3[24] ),
    .CLK(clknet_leaf_66_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[25]$_DFF_P_  (.D(\core.CPU_src1_value_a2[25] ),
    .Q(\core.CPU_src1_value_a3[25] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[26]$_DFF_P_  (.D(\core.CPU_src1_value_a2[26] ),
    .Q(\core.CPU_src1_value_a3[26] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[27]$_DFF_P_  (.D(\core.CPU_src1_value_a2[27] ),
    .Q(\core.CPU_src1_value_a3[27] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[28]$_DFF_P_  (.D(\core.CPU_src1_value_a2[28] ),
    .Q(\core.CPU_src1_value_a3[28] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[29]$_DFF_P_  (.D(\core.CPU_src1_value_a2[29] ),
    .Q(\core.CPU_src1_value_a3[29] ),
    .CLK(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[2]$_DFF_P_  (.D(\core.CPU_src1_value_a2[2] ),
    .Q(\core.CPU_src1_value_a3[2] ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[30]$_DFF_P_  (.D(\core.CPU_src1_value_a2[30] ),
    .Q(\core.CPU_src1_value_a3[30] ),
    .CLK(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[31]$_DFF_P_  (.D(\core.CPU_src1_value_a2[31] ),
    .Q(\core.CPU_src1_value_a3[31] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[3]$_DFF_P_  (.D(net350),
    .Q(\core.CPU_src1_value_a3[3] ),
    .CLK(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[4]$_DFF_P_  (.D(\core.CPU_src1_value_a2[4] ),
    .Q(\core.CPU_src1_value_a3[4] ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[5]$_DFF_P_  (.D(\core.CPU_src1_value_a2[5] ),
    .Q(\core.CPU_src1_value_a3[5] ),
    .CLK(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[6]$_DFF_P_  (.D(\core.CPU_src1_value_a2[6] ),
    .Q(\core.CPU_src1_value_a3[6] ),
    .CLK(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[7]$_DFF_P_  (.D(\core.CPU_src1_value_a2[7] ),
    .Q(\core.CPU_src1_value_a3[7] ),
    .CLK(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[8]$_DFF_P_  (.D(\core.CPU_src1_value_a2[8] ),
    .Q(\core.CPU_src1_value_a3[8] ),
    .CLK(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src1_value_a3[9]$_DFF_P_  (.D(\core.CPU_src1_value_a2[9] ),
    .Q(\core.CPU_src1_value_a3[9] ),
    .CLK(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[0]$_DFF_P_  (.D(net380),
    .Q(\core.CPU_src2_value_a3[0] ),
    .CLK(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[10]$_DFF_P_  (.D(\core.CPU_src2_value_a2[10] ),
    .Q(\core.CPU_src2_value_a3[10] ),
    .CLK(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[11]$_DFF_P_  (.D(\core.CPU_src2_value_a2[11] ),
    .Q(\core.CPU_src2_value_a3[11] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[12]$_DFF_P_  (.D(\core.CPU_src2_value_a2[12] ),
    .Q(\core.CPU_src2_value_a3[12] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[13]$_DFF_P_  (.D(net349),
    .Q(\core.CPU_src2_value_a3[13] ),
    .CLK(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[14]$_DFF_P_  (.D(\core.CPU_src2_value_a2[14] ),
    .Q(\core.CPU_src2_value_a3[14] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[15]$_DFF_P_  (.D(\core.CPU_src2_value_a2[15] ),
    .Q(\core.CPU_src2_value_a3[15] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[16]$_DFF_P_  (.D(\core.CPU_src2_value_a2[16] ),
    .Q(\core.CPU_src2_value_a3[16] ),
    .CLK(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[17]$_DFF_P_  (.D(\core.CPU_src2_value_a2[17] ),
    .Q(\core.CPU_src2_value_a3[17] ),
    .CLK(clknet_leaf_66_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[18]$_DFF_P_  (.D(\core.CPU_src2_value_a2[18] ),
    .Q(\core.CPU_src2_value_a3[18] ),
    .CLK(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[19]$_DFF_P_  (.D(\core.CPU_src2_value_a2[19] ),
    .Q(\core.CPU_src2_value_a3[19] ),
    .CLK(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[1]$_DFF_P_  (.D(\core.CPU_src2_value_a2[1] ),
    .Q(\core.CPU_src2_value_a3[1] ),
    .CLK(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[20]$_DFF_P_  (.D(\core.CPU_src2_value_a2[20] ),
    .Q(\core.CPU_src2_value_a3[20] ),
    .CLK(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[21]$_DFF_P_  (.D(\core.CPU_src2_value_a2[21] ),
    .Q(\core.CPU_src2_value_a3[21] ),
    .CLK(clknet_leaf_68_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[22]$_DFF_P_  (.D(\core.CPU_src2_value_a2[22] ),
    .Q(\core.CPU_src2_value_a3[22] ),
    .CLK(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[23]$_DFF_P_  (.D(\core.CPU_src2_value_a2[23] ),
    .Q(\core.CPU_src2_value_a3[23] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[24]$_DFF_P_  (.D(\core.CPU_src2_value_a2[24] ),
    .Q(\core.CPU_src2_value_a3[24] ),
    .CLK(clknet_leaf_66_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[25]$_DFF_P_  (.D(\core.CPU_src2_value_a2[25] ),
    .Q(\core.CPU_src2_value_a3[25] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[26]$_DFF_P_  (.D(\core.CPU_src2_value_a2[26] ),
    .Q(\core.CPU_src2_value_a3[26] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[27]$_DFF_P_  (.D(\core.CPU_src2_value_a2[27] ),
    .Q(\core.CPU_src2_value_a3[27] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[28]$_DFF_P_  (.D(\core.CPU_src2_value_a2[28] ),
    .Q(\core.CPU_src2_value_a3[28] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[29]$_DFF_P_  (.D(\core.CPU_src2_value_a2[29] ),
    .Q(\core.CPU_src2_value_a3[29] ),
    .CLK(clknet_leaf_68_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[2]$_DFF_P_  (.D(\core.CPU_src2_value_a2[2] ),
    .Q(\core.CPU_src2_value_a3[2] ),
    .CLK(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[30]$_DFF_P_  (.D(\core.CPU_src2_value_a2[30] ),
    .Q(\core.CPU_src2_value_a3[30] ),
    .CLK(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[31]$_DFF_P_  (.D(\core.CPU_src2_value_a2[31] ),
    .Q(\core.CPU_src2_value_a3[31] ),
    .CLK(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[3]$_DFF_P_  (.D(\core.CPU_src2_value_a2[3] ),
    .Q(\core.CPU_src2_value_a3[3] ),
    .CLK(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[4]$_DFF_P_  (.D(\core.CPU_src2_value_a2[4] ),
    .Q(\core.CPU_src2_value_a3[4] ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[5]$_DFF_P_  (.D(\core.CPU_src2_value_a2[5] ),
    .Q(\core.CPU_src2_value_a3[5] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[6]$_DFF_P_  (.D(\core.CPU_src2_value_a2[6] ),
    .Q(\core.CPU_src2_value_a3[6] ),
    .CLK(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[7]$_DFF_P_  (.D(\core.CPU_src2_value_a2[7] ),
    .Q(\core.CPU_src2_value_a3[7] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[8]$_DFF_P_  (.D(\core.CPU_src2_value_a2[8] ),
    .Q(\core.CPU_src2_value_a3[8] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a3[9]$_DFF_P_  (.D(\core.CPU_src2_value_a2[9] ),
    .Q(\core.CPU_src2_value_a3[9] ),
    .CLK(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[0]$_DFF_P_  (.D(\core.CPU_src2_value_a3[0] ),
    .Q(\core.CPU_dmem_wr_data_a4[0] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[10]$_DFF_P_  (.D(\core.CPU_src2_value_a3[10] ),
    .Q(\core.CPU_dmem_wr_data_a4[10] ),
    .CLK(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[11]$_DFF_P_  (.D(\core.CPU_src2_value_a3[11] ),
    .Q(\core.CPU_dmem_wr_data_a4[11] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[12]$_DFF_P_  (.D(\core.CPU_src2_value_a3[12] ),
    .Q(\core.CPU_dmem_wr_data_a4[12] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[13]$_DFF_P_  (.D(\core.CPU_src2_value_a3[13] ),
    .Q(\core.CPU_dmem_wr_data_a4[13] ),
    .CLK(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[14]$_DFF_P_  (.D(\core.CPU_src2_value_a3[14] ),
    .Q(\core.CPU_dmem_wr_data_a4[14] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[15]$_DFF_P_  (.D(\core.CPU_src2_value_a3[15] ),
    .Q(\core.CPU_dmem_wr_data_a4[15] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[16]$_DFF_P_  (.D(\core.CPU_src2_value_a3[16] ),
    .Q(\core.CPU_dmem_wr_data_a4[16] ),
    .CLK(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[17]$_DFF_P_  (.D(\core.CPU_src2_value_a3[17] ),
    .Q(\core.CPU_dmem_wr_data_a4[17] ),
    .CLK(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[18]$_DFF_P_  (.D(\core.CPU_src2_value_a3[18] ),
    .Q(\core.CPU_dmem_wr_data_a4[18] ),
    .CLK(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[19]$_DFF_P_  (.D(\core.CPU_src2_value_a3[19] ),
    .Q(\core.CPU_dmem_wr_data_a4[19] ),
    .CLK(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[1]$_DFF_P_  (.D(\core.CPU_src2_value_a3[1] ),
    .Q(\core.CPU_dmem_wr_data_a4[1] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[20]$_DFF_P_  (.D(\core.CPU_src2_value_a3[20] ),
    .Q(\core.CPU_dmem_wr_data_a4[20] ),
    .CLK(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[21]$_DFF_P_  (.D(\core.CPU_src2_value_a3[21] ),
    .Q(\core.CPU_dmem_wr_data_a4[21] ),
    .CLK(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[22]$_DFF_P_  (.D(\core.CPU_src2_value_a3[22] ),
    .Q(\core.CPU_dmem_wr_data_a4[22] ),
    .CLK(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[23]$_DFF_P_  (.D(\core.CPU_src2_value_a3[23] ),
    .Q(\core.CPU_dmem_wr_data_a4[23] ),
    .CLK(clknet_leaf_66_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[24]$_DFF_P_  (.D(\core.CPU_src2_value_a3[24] ),
    .Q(\core.CPU_dmem_wr_data_a4[24] ),
    .CLK(clknet_leaf_66_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[25]$_DFF_P_  (.D(\core.CPU_src2_value_a3[25] ),
    .Q(\core.CPU_dmem_wr_data_a4[25] ),
    .CLK(clknet_leaf_68_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[26]$_DFF_P_  (.D(\core.CPU_src2_value_a3[26] ),
    .Q(\core.CPU_dmem_wr_data_a4[26] ),
    .CLK(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[27]$_DFF_P_  (.D(\core.CPU_src2_value_a3[27] ),
    .Q(\core.CPU_dmem_wr_data_a4[27] ),
    .CLK(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[28]$_DFF_P_  (.D(\core.CPU_src2_value_a3[28] ),
    .Q(\core.CPU_dmem_wr_data_a4[28] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[29]$_DFF_P_  (.D(net586),
    .Q(\core.CPU_dmem_wr_data_a4[29] ),
    .CLK(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[2]$_DFF_P_  (.D(\core.CPU_src2_value_a3[2] ),
    .Q(\core.CPU_dmem_wr_data_a4[2] ),
    .CLK(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[30]$_DFF_P_  (.D(\core.CPU_src2_value_a3[30] ),
    .Q(\core.CPU_dmem_wr_data_a4[30] ),
    .CLK(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[31]$_DFF_P_  (.D(net585),
    .Q(\core.CPU_dmem_wr_data_a4[31] ),
    .CLK(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[3]$_DFF_P_  (.D(\core.CPU_src2_value_a3[3] ),
    .Q(\core.CPU_dmem_wr_data_a4[3] ),
    .CLK(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[4]$_DFF_P_  (.D(\core.CPU_src2_value_a3[4] ),
    .Q(\core.CPU_dmem_wr_data_a4[4] ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[5]$_DFF_P_  (.D(\core.CPU_src2_value_a3[5] ),
    .Q(\core.CPU_dmem_wr_data_a4[5] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[6]$_DFF_P_  (.D(\core.CPU_src2_value_a3[6] ),
    .Q(\core.CPU_dmem_wr_data_a4[6] ),
    .CLK(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[7]$_DFF_P_  (.D(\core.CPU_src2_value_a3[7] ),
    .Q(\core.CPU_dmem_wr_data_a4[7] ),
    .CLK(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[8]$_DFF_P_  (.D(\core.CPU_src2_value_a3[8] ),
    .Q(\core.CPU_dmem_wr_data_a4[8] ),
    .CLK(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_src2_value_a4[9]$_DFF_P_  (.D(\core.CPU_src2_value_a3[9] ),
    .Q(\core.CPU_dmem_wr_data_a4[9] ),
    .CLK(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_valid_a4$_DFF_P_  (.D(net536),
    .Q(\core.CPU_valid_a4 ),
    .CLK(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_valid_load_a4$_DFF_P_  (.D(\core.CPU_valid_load_a3 ),
    .Q(\core.CPU_dmem_rd_en_a4 ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_valid_load_a5$_DFF_P_  (.D(\core.CPU_dmem_rd_en_a4 ),
    .Q(\core.CPU_valid_load_a5 ),
    .CLK(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_valid_taken_br_a4$_DFF_P_  (.D(net377),
    .Q(\core.CPU_valid_taken_br_a4 ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.CPU_valid_taken_br_a5$_DFF_P_  (.D(\core.CPU_valid_taken_br_a4 ),
    .Q(\core.CPU_valid_taken_br_a5 ),
    .CLK(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[0]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][0] ),
    .Q(\RV_TO_DAC[0] ),
    .CLK(clknet_leaf_112_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[1]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][1] ),
    .Q(\RV_TO_DAC[1] ),
    .CLK(clknet_leaf_112_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[2]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][2] ),
    .Q(\RV_TO_DAC[2] ),
    .CLK(clknet_leaf_112_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[3]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][3] ),
    .Q(\RV_TO_DAC[3] ),
    .CLK(clknet_leaf_111_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[4]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][4] ),
    .Q(\RV_TO_DAC[4] ),
    .CLK(clknet_leaf_112_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[5]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][5] ),
    .Q(\RV_TO_DAC[5] ),
    .CLK(clknet_leaf_112_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[6]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][6] ),
    .Q(\RV_TO_DAC[6] ),
    .CLK(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[7]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][7] ),
    .Q(\RV_TO_DAC[7] ),
    .CLK(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[8]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][8] ),
    .Q(\RV_TO_DAC[8] ),
    .CLK(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__dfxtp_1 \core.OUT[9]$_DFF_P_  (.D(\core.CPU_Xreg_value_a5[17][9] ),
    .Q(\RV_TO_DAC[9] ),
    .CLK(clknet_leaf_87_CLK));
 avsddac dac (.VREFH(net8),
    .OUT(net10),
    .D({net563,
    \RV_TO_DAC[8] ,
    \RV_TO_DAC[7] ,
    \RV_TO_DAC[6] ,
    \RV_TO_DAC[5] ,
    \RV_TO_DAC[4] ,
    \RV_TO_DAC[3] ,
    \RV_TO_DAC[2] ,
    \RV_TO_DAC[1] ,
    \RV_TO_DAC[0] }));
 avsdpll pll (.ENb_CP(net4),
    .CLK(CLK),
    .ENb_VCO(net5),
    .VCO_IN(net7),
    .REF(net6));
 sky130_fd_sc_hd__conb_1 \core.CPU_is_load_a2$_DFF_P__1  (.LO(net));
 sky130_fd_sc_hd__conb_1 \core.CPU_is_s_instr_a2$_DFF_P__2  (.LO(net1));
 sky130_fd_sc_hd__conb_1 \core.CPU_is_sll_a2$_DFF_P__3  (.LO(net2));
 sky130_fd_sc_hd__conb_1 \core.CPU_is_slli_a2$_DFF_P__4  (.LO(net3));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input5 (.A(ENb_CP),
    .X(net4));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input6 (.A(ENb_VCO),
    .X(net5));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input7 (.A(REF),
    .X(net6));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input8 (.A(VCO_IN),
    .X(net7));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input9 (.A(VREFH),
    .X(net8));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input10 (.A(reset),
    .X(net9));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output11 (.A(net10),
    .X(OUT));
 sky130_fd_sc_hd__buf_4 place353 (.A(_03661_),
    .X(net352));
 sky130_fd_sc_hd__buf_4 place363 (.A(_03707_),
    .X(net362));
 sky130_fd_sc_hd__buf_4 place359 (.A(_03091_),
    .X(net358));
 sky130_fd_sc_hd__buf_4 place360 (.A(_03042_),
    .X(net359));
 sky130_fd_sc_hd__buf_4 place367 (.A(_03522_),
    .X(net366));
 sky130_fd_sc_hd__buf_4 place374 (.A(_03537_),
    .X(net373));
 sky130_fd_sc_hd__buf_4 place378 (.A(_01167_),
    .X(net377));
 sky130_fd_sc_hd__buf_4 place412 (.A(_04237_),
    .X(net411));
 sky130_fd_sc_hd__buf_4 place416 (.A(_04124_),
    .X(net415));
 sky130_fd_sc_hd__buf_4 place414 (.A(_04181_),
    .X(net413));
 sky130_fd_sc_hd__buf_4 place415 (.A(_04127_),
    .X(net414));
 sky130_fd_sc_hd__buf_4 place417 (.A(_04080_),
    .X(net416));
 sky130_fd_sc_hd__buf_4 place419 (.A(_04021_),
    .X(net418));
 sky130_fd_sc_hd__buf_4 place422 (.A(_03955_),
    .X(net421));
 sky130_fd_sc_hd__buf_4 place423 (.A(_03901_),
    .X(net422));
 sky130_fd_sc_hd__buf_4 place427 (.A(_03751_),
    .X(net426));
 sky130_fd_sc_hd__buf_4 place432 (.A(net430),
    .X(net431));
 sky130_fd_sc_hd__buf_4 place428 (.A(_02859_),
    .X(net427));
 sky130_fd_sc_hd__buf_4 place433 (.A(_04399_),
    .X(net432));
 sky130_fd_sc_hd__buf_4 place437 (.A(_03435_),
    .X(net436));
 sky130_fd_sc_hd__buf_4 place442 (.A(_02530_),
    .X(net441));
 sky130_fd_sc_hd__buf_4 place436 (.A(_02665_),
    .X(net435));
 sky130_fd_sc_hd__buf_4 place438 (.A(_03230_),
    .X(net437));
 sky130_fd_sc_hd__buf_4 place439 (.A(_03048_),
    .X(net438));
 sky130_fd_sc_hd__buf_4 place443 (.A(_02430_),
    .X(net442));
 sky130_fd_sc_hd__buf_4 place440 (.A(_02814_),
    .X(net439));
 sky130_fd_sc_hd__buf_4 place441 (.A(_02544_),
    .X(net440));
 sky130_fd_sc_hd__buf_4 place445 (.A(_02277_),
    .X(net444));
 sky130_fd_sc_hd__buf_4 place446 (.A(_02202_),
    .X(net445));
 sky130_fd_sc_hd__buf_4 place447 (.A(_02123_),
    .X(net446));
 sky130_fd_sc_hd__buf_4 place448 (.A(_02050_),
    .X(net447));
 sky130_fd_sc_hd__buf_4 place449 (.A(_01967_),
    .X(net448));
 sky130_fd_sc_hd__buf_4 place450 (.A(_01893_),
    .X(net449));
 sky130_fd_sc_hd__buf_4 place451 (.A(_01813_),
    .X(net450));
 sky130_fd_sc_hd__buf_4 place452 (.A(_01735_),
    .X(net451));
 sky130_fd_sc_hd__buf_4 place453 (.A(_01661_),
    .X(net452));
 sky130_fd_sc_hd__buf_4 place454 (.A(_01583_),
    .X(net453));
 sky130_fd_sc_hd__buf_4 place455 (.A(_01508_),
    .X(net454));
 sky130_fd_sc_hd__buf_4 place456 (.A(_01427_),
    .X(net455));
 sky130_fd_sc_hd__buf_4 place457 (.A(_01352_),
    .X(net456));
 sky130_fd_sc_hd__buf_4 place458 (.A(_01200_),
    .X(net457));
 sky130_fd_sc_hd__buf_4 place459 (.A(_04884_),
    .X(net458));
 sky130_fd_sc_hd__buf_4 place463 (.A(_04752_),
    .X(net462));
 sky130_fd_sc_hd__buf_4 place485 (.A(_02355_),
    .X(net484));
 sky130_fd_sc_hd__buf_4 place466 (.A(_04492_),
    .X(net465));
 sky130_fd_sc_hd__buf_4 place465 (.A(_04521_),
    .X(net464));
 sky130_fd_sc_hd__buf_4 place487 (.A(_02352_),
    .X(net486));
 sky130_fd_sc_hd__buf_4 place462 (.A(_04760_),
    .X(net461));
 sky130_fd_sc_hd__buf_4 place460 (.A(_04816_),
    .X(net459));
 sky130_fd_sc_hd__buf_4 place489 (.A(_02280_),
    .X(net488));
 sky130_fd_sc_hd__buf_4 place461 (.A(_04791_),
    .X(net460));
 sky130_fd_sc_hd__buf_4 place491 (.A(_02275_),
    .X(net490));
 sky130_fd_sc_hd__buf_4 place435 (.A(_04399_),
    .X(net434));
 sky130_fd_sc_hd__buf_4 place434 (.A(net432),
    .X(net433));
 sky130_fd_sc_hd__buf_4 place408 (.A(_04490_),
    .X(net407));
 sky130_fd_sc_hd__buf_4 place492 (.A(_02201_),
    .X(net491));
 sky130_fd_sc_hd__buf_4 place406 (.A(_04533_),
    .X(net405));
 sky130_fd_sc_hd__buf_4 place403 (.A(_04588_),
    .X(net402));
 sky130_fd_sc_hd__buf_4 place494 (.A(_02198_),
    .X(net493));
 sky130_fd_sc_hd__buf_4 place496 (.A(_02126_),
    .X(net495));
 sky130_fd_sc_hd__buf_4 place498 (.A(_02122_),
    .X(net497));
 sky130_fd_sc_hd__buf_4 place402 (.A(_04678_),
    .X(net401));
 sky130_fd_sc_hd__buf_4 place401 (.A(_04697_),
    .X(net400));
 sky130_fd_sc_hd__buf_4 place400 (.A(_04723_),
    .X(net399));
 sky130_fd_sc_hd__buf_4 place500 (.A(_02049_),
    .X(net499));
 sky130_fd_sc_hd__buf_4 place399 (.A(_04732_),
    .X(net398));
 sky130_fd_sc_hd__buf_4 place502 (.A(_02046_),
    .X(net501));
 sky130_fd_sc_hd__buf_4 place398 (.A(_04871_),
    .X(net397));
 sky130_fd_sc_hd__buf_4 place397 (.A(_04880_),
    .X(net396));
 sky130_fd_sc_hd__buf_4 place504 (.A(_01970_),
    .X(net503));
 sky130_fd_sc_hd__buf_4 place506 (.A(_01965_),
    .X(net505));
 sky130_fd_sc_hd__buf_4 place390 (.A(_04240_),
    .X(net389));
 sky130_fd_sc_hd__buf_4 place389 (.A(_04514_),
    .X(net388));
 sky130_fd_sc_hd__buf_4 place387 (.A(_04717_),
    .X(net386));
 sky130_fd_sc_hd__buf_4 place385 (.A(_04992_),
    .X(net384));
 sky130_fd_sc_hd__buf_4 place381 (.A(\core.CPU_src2_value_a2[0] ),
    .X(net380));
 sky130_fd_sc_hd__buf_4 place508 (.A(_01891_),
    .X(net507));
 sky130_fd_sc_hd__buf_4 place384 (.A(_05015_),
    .X(net383));
 sky130_fd_sc_hd__buf_4 place386 (.A(_04981_),
    .X(net385));
 sky130_fd_sc_hd__buf_4 place352 (.A(_03725_),
    .X(net351));
 sky130_fd_sc_hd__buf_4 place510 (.A(_01888_),
    .X(net509));
 sky130_fd_sc_hd__buf_4 place369 (.A(_03276_),
    .X(net368));
 sky130_fd_sc_hd__buf_4 place512 (.A(_01816_),
    .X(net511));
 sky130_fd_sc_hd__buf_4 place345 (.A(_03696_),
    .X(net344));
 sky130_fd_sc_hd__buf_4 place351 (.A(\core.CPU_src1_value_a2[3] ),
    .X(net350));
 sky130_fd_sc_hd__buf_4 place515 (.A(_01811_),
    .X(net514));
 sky130_fd_sc_hd__buf_4 place410 (.A(_04298_),
    .X(net409));
 sky130_fd_sc_hd__buf_4 place514 (.A(_01811_),
    .X(net513));
 sky130_fd_sc_hd__buf_4 place388 (.A(_04656_),
    .X(net387));
 sky130_fd_sc_hd__buf_4 place405 (.A(_04553_),
    .X(net404));
 sky130_fd_sc_hd__buf_4 place617 (.A(\core.CPU_Xreg_value_a4[17][5] ),
    .X(net616));
 sky130_fd_sc_hd__buf_4 place516 (.A(_01738_),
    .X(net515));
 sky130_fd_sc_hd__buf_4 place350 (.A(\core.CPU_src2_value_a2[13] ),
    .X(net349));
 sky130_fd_sc_hd__buf_4 place383 (.A(_05025_),
    .X(net382));
 sky130_fd_sc_hd__buf_4 place382 (.A(_04570_),
    .X(net381));
 sky130_fd_sc_hd__buf_4 place518 (.A(_01734_),
    .X(net517));
 sky130_fd_sc_hd__buf_4 place619 (.A(\core.CPU_Xreg_value_a4[17][2] ),
    .X(net618));
 sky130_fd_sc_hd__buf_4 place618 (.A(\core.CPU_Xreg_value_a4[17][4] ),
    .X(net617));
 sky130_fd_sc_hd__buf_4 place519 (.A(_01660_),
    .X(net518));
 sky130_fd_sc_hd__buf_4 place620 (.A(\core.CPU_Xreg_value_a4[17][1] ),
    .X(net619));
 sky130_fd_sc_hd__buf_4 place621 (.A(\core.CPU_Xreg_value_a4[17][0] ),
    .X(net620));
 sky130_fd_sc_hd__buf_4 place520 (.A(_01657_),
    .X(net519));
 sky130_fd_sc_hd__buf_4 place522 (.A(_01586_),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_CLK (.A(clknet_4_12_0_CLK),
    .X(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__buf_4 place523 (.A(_01582_),
    .X(net522));
 sky130_fd_sc_hd__buf_4 place616 (.A(\core.CPU_imem_rd_addr_a1[2] ),
    .X(net615));
 sky130_fd_sc_hd__buf_4 place615 (.A(\core.CPU_imem_rd_addr_a1[3] ),
    .X(net614));
 sky130_fd_sc_hd__buf_4 place524 (.A(_01507_),
    .X(net523));
 sky130_fd_sc_hd__buf_4 place607 (.A(\core.CPU_reset_a3 ),
    .X(net606));
 sky130_fd_sc_hd__buf_4 place526 (.A(_01504_),
    .X(net525));
 sky130_fd_sc_hd__buf_4 place527 (.A(_01430_),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_CLK (.A(clknet_4_13_0_CLK),
    .X(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__buf_12 place608 (.A(net606),
    .X(net607));
 sky130_fd_sc_hd__buf_4 place550 (.A(_02644_),
    .X(net549));
 sky130_fd_sc_hd__buf_4 place528 (.A(_01426_),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_CLK (.A(clknet_4_12_0_CLK),
    .X(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__buf_4 place554 (.A(_02578_),
    .X(net553));
 sky130_fd_sc_hd__buf_4 place558 (.A(_02512_),
    .X(net557));
 sky130_fd_sc_hd__buf_4 place548 (.A(_02791_),
    .X(net547));
 sky130_fd_sc_hd__buf_4 place530 (.A(_01351_),
    .X(net529));
 sky130_fd_sc_hd__buf_4 place547 (.A(_02819_),
    .X(net546));
 sky130_fd_sc_hd__buf_4 place532 (.A(_01348_),
    .X(net531));
 sky130_fd_sc_hd__buf_4 place534 (.A(_01207_),
    .X(net533));
 sky130_fd_sc_hd__buf_4 place545 (.A(_04406_),
    .X(net544));
 sky130_fd_sc_hd__buf_4 place535 (.A(_01199_),
    .X(net534));
 sky130_fd_sc_hd__buf_4 place544 (.A(_04410_),
    .X(net543));
 sky130_fd_sc_hd__buf_4 place536 (.A(_01115_),
    .X(net535));
 sky130_fd_sc_hd__buf_4 place538 (.A(_04804_),
    .X(net537));
 sky130_fd_sc_hd__buf_4 place539 (.A(_04759_),
    .X(net538));
 sky130_fd_sc_hd__buf_4 place557 (.A(_02536_),
    .X(net556));
 sky130_fd_sc_hd__buf_4 place555 (.A(_02570_),
    .X(net554));
 sky130_fd_sc_hd__buf_4 place556 (.A(_02537_),
    .X(net555));
 sky130_fd_sc_hd__buf_4 place561 (.A(_01203_),
    .X(net560));
 sky130_fd_sc_hd__buf_4 place563 (.A(_01114_),
    .X(net562));
 sky130_fd_sc_hd__buf_4 place562 (.A(_01191_),
    .X(net561));
 sky130_fd_sc_hd__buf_4 place598 (.A(\core.CPU_rf_rd_index1_a2[0] ),
    .X(net597));
 sky130_fd_sc_hd__buf_4 place564 (.A(\RV_TO_DAC[9] ),
    .X(net563));
 sky130_fd_sc_hd__buf_4 place590 (.A(\core.CPU_rf_rd_index2_a2[1] ),
    .X(net589));
 sky130_fd_sc_hd__buf_4 place592 (.A(\core.CPU_rf_rd_index2_a2[0] ),
    .X(net591));
 sky130_fd_sc_hd__buf_4 place594 (.A(\core.CPU_rf_rd_index1_a2[4] ),
    .X(net593));
 sky130_fd_sc_hd__buf_4 place596 (.A(\core.CPU_rf_rd_index1_a2[1] ),
    .X(net595));
 sky130_fd_sc_hd__buf_4 place599 (.A(\core.CPU_rf_rd_index1_a2[0] ),
    .X(net598));
 sky130_fd_sc_hd__buf_4 place601 (.A(\core.CPU_reset_a4 ),
    .X(net600));
 sky130_fd_sc_hd__buf_4 place600 (.A(\core.CPU_reset_a4 ),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_CLK (.A(clknet_4_12_0_CLK),
    .X(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__buf_4 place614 (.A(\core.CPU_imm_a3[12] ),
    .X(net613));
 sky130_fd_sc_hd__buf_4 place610 (.A(\core.CPU_is_sub_a3 ),
    .X(net609));
 sky130_fd_sc_hd__buf_4 place609 (.A(\core.CPU_reset_a1 ),
    .X(net608));
 sky130_fd_sc_hd__buf_4 place613 (.A(\core.CPU_is_add_a3 ),
    .X(net612));
 sky130_fd_sc_hd__buf_4 place611 (.A(\core.CPU_is_slli_a3 ),
    .X(net610));
 sky130_fd_sc_hd__buf_4 place612 (.A(\core.CPU_is_addi_a3 ),
    .X(net611));
 sky130_fd_sc_hd__buf_4 place346 (.A(_03580_),
    .X(net345));
 sky130_fd_sc_hd__buf_4 place347 (.A(_02957_),
    .X(net346));
 sky130_fd_sc_hd__buf_4 place348 (.A(_02868_),
    .X(net347));
 sky130_fd_sc_hd__buf_4 place349 (.A(_02642_),
    .X(net348));
 sky130_fd_sc_hd__buf_4 place354 (.A(_03420_),
    .X(net353));
 sky130_fd_sc_hd__buf_4 place355 (.A(_03353_),
    .X(net354));
 sky130_fd_sc_hd__buf_4 place356 (.A(_03231_),
    .X(net355));
 sky130_fd_sc_hd__buf_4 place357 (.A(_03191_),
    .X(net356));
 sky130_fd_sc_hd__buf_4 place358 (.A(_03143_),
    .X(net357));
 sky130_fd_sc_hd__buf_4 place361 (.A(_02767_),
    .X(net360));
 sky130_fd_sc_hd__buf_4 place362 (.A(_02719_),
    .X(net361));
 sky130_fd_sc_hd__buf_4 place364 (.A(_03642_),
    .X(net363));
 sky130_fd_sc_hd__buf_4 place365 (.A(_03625_),
    .X(net364));
 sky130_fd_sc_hd__buf_4 place366 (.A(_03610_),
    .X(net365));
 sky130_fd_sc_hd__buf_4 place368 (.A(_03407_),
    .X(net367));
 sky130_fd_sc_hd__buf_4 place370 (.A(_03229_),
    .X(net369));
 sky130_fd_sc_hd__buf_4 place372 (.A(_03677_),
    .X(net371));
 sky130_fd_sc_hd__buf_4 place371 (.A(_02760_),
    .X(net370));
 sky130_fd_sc_hd__buf_4 place373 (.A(\core.CPU_result_a3[3] ),
    .X(net372));
 sky130_fd_sc_hd__buf_4 place380 (.A(_04808_),
    .X(net379));
 sky130_fd_sc_hd__buf_4 place375 (.A(\core.CPU_src1_value_a2[0] ),
    .X(net374));
 sky130_fd_sc_hd__buf_4 place376 (.A(_03100_),
    .X(net375));
 sky130_fd_sc_hd__buf_4 place377 (.A(_03074_),
    .X(net376));
 sky130_fd_sc_hd__buf_4 place379 (.A(_04863_),
    .X(net378));
 sky130_fd_sc_hd__buf_4 place391 (.A(_03836_),
    .X(net390));
 sky130_fd_sc_hd__buf_4 place395 (.A(_02543_),
    .X(net394));
 sky130_fd_sc_hd__buf_4 place392 (.A(_03471_),
    .X(net391));
 sky130_fd_sc_hd__buf_4 place393 (.A(_03177_),
    .X(net392));
 sky130_fd_sc_hd__buf_4 place394 (.A(_03109_),
    .X(net393));
 sky130_fd_sc_hd__buf_4 place396 (.A(_04999_),
    .X(net395));
 sky130_fd_sc_hd__buf_4 place404 (.A(_04560_),
    .X(net403));
 sky130_fd_sc_hd__buf_4 place407 (.A(_04498_),
    .X(net406));
 sky130_fd_sc_hd__buf_4 place409 (.A(_04460_),
    .X(net408));
 sky130_fd_sc_hd__buf_4 place411 (.A(_04290_),
    .X(net410));
 sky130_fd_sc_hd__buf_4 place413 (.A(_04188_),
    .X(net412));
 sky130_fd_sc_hd__buf_4 place418 (.A(_04071_),
    .X(net417));
 sky130_fd_sc_hd__buf_4 place420 (.A(_04018_),
    .X(net419));
 sky130_fd_sc_hd__buf_4 place421 (.A(_03963_),
    .X(net420));
 sky130_fd_sc_hd__buf_4 place424 (.A(_03893_),
    .X(net423));
 sky130_fd_sc_hd__buf_4 place425 (.A(_03831_),
    .X(net424));
 sky130_fd_sc_hd__buf_4 place426 (.A(_03761_),
    .X(net425));
 sky130_fd_sc_hd__buf_4 place429 (.A(_02563_),
    .X(net428));
 sky130_fd_sc_hd__buf_4 place430 (.A(_02558_),
    .X(net429));
 sky130_fd_sc_hd__buf_4 place431 (.A(_04745_),
    .X(net430));
 sky130_fd_sc_hd__buf_4 place444 (.A(_02356_),
    .X(net443));
 sky130_fd_sc_hd__buf_4 place464 (.A(_04737_),
    .X(net463));
 sky130_fd_sc_hd__buf_4 place468 (.A(_04442_),
    .X(net467));
 sky130_fd_sc_hd__buf_4 place472 (.A(_04416_),
    .X(net471));
 sky130_fd_sc_hd__buf_4 place475 (.A(_02919_),
    .X(net474));
 sky130_fd_sc_hd__buf_4 place474 (.A(_02931_),
    .X(net473));
 sky130_fd_sc_hd__buf_4 place476 (.A(_02917_),
    .X(net475));
 sky130_fd_sc_hd__buf_4 place477 (.A(_02864_),
    .X(net476));
 sky130_fd_sc_hd__buf_4 place478 (.A(_02681_),
    .X(net477));
 sky130_fd_sc_hd__buf_4 place480 (.A(_02533_),
    .X(net479));
 sky130_fd_sc_hd__buf_4 place482 (.A(_02521_),
    .X(net481));
 sky130_fd_sc_hd__buf_4 place483 (.A(_02433_),
    .X(net482));
 sky130_fd_sc_hd__buf_4 place486 (.A(_02355_),
    .X(net485));
 sky130_fd_sc_hd__buf_4 place484 (.A(_02428_),
    .X(net483));
 sky130_fd_sc_hd__buf_4 place467 (.A(_04472_),
    .X(net466));
 sky130_fd_sc_hd__buf_4 place469 (.A(_04439_),
    .X(net468));
 sky130_fd_sc_hd__buf_4 place470 (.A(_04429_),
    .X(net469));
 sky130_fd_sc_hd__buf_4 place471 (.A(_04429_),
    .X(net470));
 sky130_fd_sc_hd__buf_4 place473 (.A(_04411_),
    .X(net472));
 sky130_fd_sc_hd__buf_4 place479 (.A(_02587_),
    .X(net478));
 sky130_fd_sc_hd__buf_4 place481 (.A(_02528_),
    .X(net480));
 sky130_fd_sc_hd__buf_4 place488 (.A(_02352_),
    .X(net487));
 sky130_fd_sc_hd__buf_4 place490 (.A(net488),
    .X(net489));
 sky130_fd_sc_hd__buf_4 place493 (.A(net491),
    .X(net492));
 sky130_fd_sc_hd__buf_4 place495 (.A(net493),
    .X(net494));
 sky130_fd_sc_hd__buf_4 place497 (.A(_02126_),
    .X(net496));
 sky130_fd_sc_hd__buf_4 place499 (.A(net497),
    .X(net498));
 sky130_fd_sc_hd__buf_4 place501 (.A(net499),
    .X(net500));
 sky130_fd_sc_hd__buf_4 place503 (.A(net501),
    .X(net502));
 sky130_fd_sc_hd__buf_4 place505 (.A(net503),
    .X(net504));
 sky130_fd_sc_hd__buf_4 place507 (.A(net505),
    .X(net506));
 sky130_fd_sc_hd__buf_4 place509 (.A(net507),
    .X(net508));
 sky130_fd_sc_hd__buf_4 place511 (.A(net509),
    .X(net510));
 sky130_fd_sc_hd__buf_4 place513 (.A(_01816_),
    .X(net512));
 sky130_fd_sc_hd__buf_4 place517 (.A(net515),
    .X(net516));
 sky130_fd_sc_hd__buf_4 place521 (.A(net519),
    .X(net520));
 sky130_fd_sc_hd__buf_4 place525 (.A(net523),
    .X(net524));
 sky130_fd_sc_hd__buf_4 place529 (.A(net527),
    .X(net528));
 sky130_fd_sc_hd__buf_4 place531 (.A(net529),
    .X(net530));
 sky130_fd_sc_hd__buf_4 place533 (.A(net531),
    .X(net532));
 sky130_fd_sc_hd__buf_4 place537 (.A(net535),
    .X(net536));
 sky130_fd_sc_hd__buf_4 place540 (.A(_04751_),
    .X(net539));
 sky130_fd_sc_hd__buf_4 place541 (.A(_04748_),
    .X(net540));
 sky130_fd_sc_hd__buf_4 place542 (.A(_04436_),
    .X(net541));
 sky130_fd_sc_hd__buf_4 place543 (.A(_04419_),
    .X(net542));
 sky130_fd_sc_hd__buf_4 place546 (.A(net544),
    .X(net545));
 sky130_fd_sc_hd__buf_4 place549 (.A(_02671_),
    .X(net548));
 sky130_fd_sc_hd__buf_4 place551 (.A(net549),
    .X(net550));
 sky130_fd_sc_hd__buf_4 place552 (.A(_02644_),
    .X(net551));
 sky130_fd_sc_hd__buf_4 place553 (.A(net551),
    .X(net552));
 sky130_fd_sc_hd__buf_4 place559 (.A(_01206_),
    .X(net558));
 sky130_fd_sc_hd__buf_4 place560 (.A(net558),
    .X(net559));
 sky130_fd_sc_hd__buf_4 place565 (.A(\core.CPU_dmem_wr_data_a4[9] ),
    .X(net564));
 sky130_fd_sc_hd__buf_4 place566 (.A(\core.CPU_dmem_wr_data_a4[8] ),
    .X(net565));
 sky130_fd_sc_hd__buf_4 place567 (.A(\core.CPU_dmem_wr_data_a4[7] ),
    .X(net566));
 sky130_fd_sc_hd__buf_4 place568 (.A(\core.CPU_dmem_wr_data_a4[6] ),
    .X(net567));
 sky130_fd_sc_hd__buf_4 place569 (.A(\core.CPU_dmem_wr_data_a4[2] ),
    .X(net568));
 sky130_fd_sc_hd__buf_4 place570 (.A(\core.CPU_dmem_wr_data_a4[27] ),
    .X(net569));
 sky130_fd_sc_hd__buf_4 place571 (.A(\core.CPU_dmem_wr_data_a4[26] ),
    .X(net570));
 sky130_fd_sc_hd__buf_4 place572 (.A(\core.CPU_dmem_wr_data_a4[25] ),
    .X(net571));
 sky130_fd_sc_hd__buf_4 place573 (.A(\core.CPU_dmem_wr_data_a4[24] ),
    .X(net572));
 sky130_fd_sc_hd__buf_4 place574 (.A(\core.CPU_dmem_wr_data_a4[23] ),
    .X(net573));
 sky130_fd_sc_hd__buf_4 place575 (.A(\core.CPU_dmem_wr_data_a4[22] ),
    .X(net574));
 sky130_fd_sc_hd__buf_4 place576 (.A(\core.CPU_dmem_wr_data_a4[21] ),
    .X(net575));
 sky130_fd_sc_hd__buf_4 place577 (.A(\core.CPU_dmem_wr_data_a4[20] ),
    .X(net576));
 sky130_fd_sc_hd__buf_4 place578 (.A(\core.CPU_dmem_wr_data_a4[1] ),
    .X(net577));
 sky130_fd_sc_hd__buf_4 place579 (.A(\core.CPU_dmem_wr_data_a4[19] ),
    .X(net578));
 sky130_fd_sc_hd__buf_4 place580 (.A(\core.CPU_dmem_wr_data_a4[17] ),
    .X(net579));
 sky130_fd_sc_hd__buf_4 place581 (.A(\core.CPU_dmem_wr_data_a4[15] ),
    .X(net580));
 sky130_fd_sc_hd__buf_4 place582 (.A(\core.CPU_dmem_wr_data_a4[14] ),
    .X(net581));
 sky130_fd_sc_hd__buf_4 place583 (.A(\core.CPU_dmem_wr_data_a4[12] ),
    .X(net582));
 sky130_fd_sc_hd__buf_4 place584 (.A(\core.CPU_dmem_wr_data_a4[11] ),
    .X(net583));
 sky130_fd_sc_hd__buf_4 place585 (.A(\core.CPU_dmem_wr_data_a4[10] ),
    .X(net584));
 sky130_fd_sc_hd__buf_4 place586 (.A(\core.CPU_src2_value_a3[31] ),
    .X(net585));
 sky130_fd_sc_hd__buf_4 place587 (.A(\core.CPU_src2_value_a3[29] ),
    .X(net586));
 sky130_fd_sc_hd__buf_4 place588 (.A(\core.CPU_rf_rd_index2_a2[3] ),
    .X(net587));
 sky130_fd_sc_hd__buf_4 place589 (.A(\core.CPU_rf_rd_index2_a2[3] ),
    .X(net588));
 sky130_fd_sc_hd__buf_4 place591 (.A(\core.CPU_rf_rd_index2_a2[1] ),
    .X(net590));
 sky130_fd_sc_hd__buf_4 place593 (.A(\core.CPU_rf_rd_index2_a2[0] ),
    .X(net592));
 sky130_fd_sc_hd__buf_4 place595 (.A(net593),
    .X(net594));
 sky130_fd_sc_hd__buf_4 place597 (.A(net595),
    .X(net596));
 sky130_fd_sc_hd__buf_12 place602 (.A(net600),
    .X(net601));
 sky130_fd_sc_hd__buf_4 place603 (.A(net600),
    .X(net602));
 sky130_fd_sc_hd__buf_4 place604 (.A(\core.CPU_reset_a4 ),
    .X(net603));
 sky130_fd_sc_hd__buf_4 place605 (.A(net603),
    .X(net604));
 sky130_fd_sc_hd__buf_4 place606 (.A(net604),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_CLK (.A(clknet_4_13_0_CLK),
    .X(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_CLK (.A(clknet_4_13_0_CLK),
    .X(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_CLK (.A(clknet_4_12_0_CLK),
    .X(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_CLK (.A(clknet_4_13_0_CLK),
    .X(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_CLK (.A(clknet_4_13_0_CLK),
    .X(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_CLK (.A(clknet_4_13_0_CLK),
    .X(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_CLK (.A(clknet_4_13_0_CLK),
    .X(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_CLK (.A(clknet_4_13_0_CLK),
    .X(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_CLK (.A(clknet_4_14_0_CLK),
    .X(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_CLK (.A(clknet_4_14_0_CLK),
    .X(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_CLK (.A(clknet_4_14_0_CLK),
    .X(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_CLK (.A(clknet_4_13_0_CLK),
    .X(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_CLK (.A(clknet_4_15_0_CLK),
    .X(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_CLK (.A(clknet_4_12_0_CLK),
    .X(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_CLK (.A(clknet_4_14_0_CLK),
    .X(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_CLK (.A(clknet_4_14_0_CLK),
    .X(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_CLK (.A(clknet_4_11_0_CLK),
    .X(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_CLK (.A(clknet_4_11_0_CLK),
    .X(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_CLK (.A(clknet_4_11_0_CLK),
    .X(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_CLK (.A(clknet_4_14_0_CLK),
    .X(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_CLK (.A(clknet_4_14_0_CLK),
    .X(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_CLK (.A(clknet_4_14_0_CLK),
    .X(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_CLK (.A(clknet_4_14_0_CLK),
    .X(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_CLK (.A(clknet_4_10_0_CLK),
    .X(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_CLK (.A(clknet_4_10_0_CLK),
    .X(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_CLK (.A(clknet_4_10_0_CLK),
    .X(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_CLK (.A(clknet_4_10_0_CLK),
    .X(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_CLK (.A(clknet_4_10_0_CLK),
    .X(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_CLK (.A(clknet_4_10_0_CLK),
    .X(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_CLK (.A(clknet_4_10_0_CLK),
    .X(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_CLK (.A(clknet_4_11_0_CLK),
    .X(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_CLK (.A(clknet_4_11_0_CLK),
    .X(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_CLK (.A(clknet_4_9_0_CLK),
    .X(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_CLK (.A(clknet_4_8_0_CLK),
    .X(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_CLK (.A(clknet_4_8_0_CLK),
    .X(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_CLK (.A(clknet_4_8_0_CLK),
    .X(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_CLK (.A(clknet_4_8_0_CLK),
    .X(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_CLK (.A(clknet_4_11_0_CLK),
    .X(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_CLK (.A(clknet_4_11_0_CLK),
    .X(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_CLK (.A(clknet_4_8_0_CLK),
    .X(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_CLK (.A(clknet_4_12_0_CLK),
    .X(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_CLK (.A(clknet_4_3_0_CLK),
    .X(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_CLK (.A(clknet_4_3_0_CLK),
    .X(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_CLK (.A(clknet_4_3_0_CLK),
    .X(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_CLK (.A(clknet_4_8_0_CLK),
    .X(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_CLK (.A(clknet_4_9_0_CLK),
    .X(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_CLK (.A(clknet_4_9_0_CLK),
    .X(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_CLK (.A(clknet_4_9_0_CLK),
    .X(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_CLK (.A(clknet_4_10_0_CLK),
    .X(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_CLK (.A(clknet_4_1_0_CLK),
    .X(clknet_leaf_65_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_CLK (.A(clknet_4_1_0_CLK),
    .X(clknet_leaf_66_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_CLK (.A(clknet_4_1_0_CLK),
    .X(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_CLK (.A(clknet_4_1_0_CLK),
    .X(clknet_leaf_68_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_CLK (.A(clknet_4_3_0_CLK),
    .X(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_CLK (.A(clknet_4_0_0_CLK),
    .X(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_CLK (.A(clknet_4_2_0_CLK),
    .X(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_CLK (.A(clknet_4_2_0_CLK),
    .X(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_CLK (.A(clknet_4_0_0_CLK),
    .X(clknet_leaf_73_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_CLK (.A(clknet_4_0_0_CLK),
    .X(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_CLK (.A(clknet_4_2_0_CLK),
    .X(clknet_leaf_75_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_CLK (.A(clknet_4_0_0_CLK),
    .X(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_80_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_CLK (.A(clknet_4_0_0_CLK),
    .X(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_CLK (.A(clknet_4_2_0_CLK),
    .X(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_CLK (.A(clknet_4_6_0_CLK),
    .X(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_CLK (.A(clknet_4_6_0_CLK),
    .X(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_CLK (.A(clknet_4_7_0_CLK),
    .X(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_CLK (.A(clknet_4_2_0_CLK),
    .X(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_CLK (.A(clknet_4_3_0_CLK),
    .X(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_CLK (.A(clknet_4_3_0_CLK),
    .X(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_CLK (.A(clknet_4_3_0_CLK),
    .X(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_CLK (.A(clknet_4_6_0_CLK),
    .X(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_CLK (.A(clknet_4_6_0_CLK),
    .X(clknet_leaf_96_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_CLK (.A(clknet_4_6_0_CLK),
    .X(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_CLK (.A(clknet_4_6_0_CLK),
    .X(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_CLK (.A(clknet_4_6_0_CLK),
    .X(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_CLK (.A(clknet_4_6_0_CLK),
    .X(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_CLK (.A(clknet_4_5_0_CLK),
    .X(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_CLK (.A(clknet_4_5_0_CLK),
    .X(clknet_leaf_102_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_CLK (.A(clknet_4_5_0_CLK),
    .X(clknet_leaf_103_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_CLK (.A(clknet_4_5_0_CLK),
    .X(clknet_leaf_104_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_CLK (.A(clknet_4_5_0_CLK),
    .X(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_CLK (.A(clknet_4_4_0_CLK),
    .X(clknet_leaf_106_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_CLK (.A(clknet_4_4_0_CLK),
    .X(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_CLK (.A(clknet_4_4_0_CLK),
    .X(clknet_leaf_108_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_CLK (.A(clknet_4_5_0_CLK),
    .X(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_CLK (.A(clknet_4_4_0_CLK),
    .X(clknet_leaf_110_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_CLK (.A(clknet_4_4_0_CLK),
    .X(clknet_leaf_111_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_CLK (.A(clknet_4_4_0_CLK),
    .X(clknet_leaf_112_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (.A(CLK),
    .X(clknet_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_0_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_1_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_2_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_3_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_4_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_5_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_6_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_7_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_8_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_9_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_10_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_11_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_12_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_13_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_14_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_CLK (.A(clknet_0_CLK),
    .X(clknet_4_15_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload0 (.A(clknet_4_0_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload1 (.A(clknet_4_1_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload2 (.A(clknet_4_2_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload3 (.A(clknet_4_3_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload4 (.A(clknet_4_4_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload5 (.A(clknet_4_5_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload6 (.A(clknet_4_6_0_CLK));
 sky130_fd_sc_hd__clkinv_8 clkload7 (.A(clknet_4_7_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload8 (.A(clknet_4_8_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload9 (.A(clknet_4_9_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload10 (.A(clknet_4_10_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload11 (.A(clknet_4_11_0_CLK));
 sky130_fd_sc_hd__clkinv_16 clkload12 (.A(clknet_4_12_0_CLK));
 sky130_fd_sc_hd__inv_16 clkload13 (.A(clknet_4_13_0_CLK));
 sky130_fd_sc_hd__inv_16 clkload14 (.A(clknet_4_14_0_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload15 (.A(clknet_leaf_70_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload16 (.A(clknet_leaf_74_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload17 (.A(clknet_leaf_76_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload18 (.A(clknet_leaf_81_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload19 (.A(clknet_leaf_66_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload20 (.A(clknet_leaf_67_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload21 (.A(clknet_leaf_68_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload22 (.A(clknet_leaf_71_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload23 (.A(clknet_leaf_72_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload24 (.A(clknet_leaf_86_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload25 (.A(clknet_leaf_91_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload26 (.A(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload27 (.A(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload28 (.A(clknet_leaf_69_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload29 (.A(clknet_leaf_92_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload30 (.A(clknet_leaf_93_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload31 (.A(clknet_leaf_94_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload32 (.A(clknet_leaf_107_CLK));
 sky130_fd_sc_hd__inv_6 clkload33 (.A(clknet_leaf_110_CLK));
 sky130_fd_sc_hd__inv_6 clkload34 (.A(clknet_leaf_111_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload35 (.A(clknet_leaf_112_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload36 (.A(clknet_leaf_101_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload37 (.A(clknet_leaf_105_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload38 (.A(clknet_leaf_109_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload39 (.A(clknet_leaf_87_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload40 (.A(clknet_leaf_88_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload41 (.A(clknet_leaf_95_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload42 (.A(clknet_leaf_97_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload43 (.A(clknet_leaf_98_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload44 (.A(clknet_leaf_99_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload45 (.A(clknet_leaf_100_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload46 (.A(clknet_leaf_77_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload47 (.A(clknet_leaf_78_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload48 (.A(clknet_leaf_79_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload49 (.A(clknet_leaf_82_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload50 (.A(clknet_leaf_83_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload51 (.A(clknet_leaf_84_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload52 (.A(clknet_leaf_85_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload53 (.A(clknet_leaf_89_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload54 (.A(clknet_leaf_90_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload55 (.A(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload56 (.A(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload57 (.A(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload58 (.A(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload59 (.A(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload60 (.A(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload61 (.A(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload62 (.A(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload63 (.A(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload64 (.A(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload65 (.A(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload66 (.A(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload67 (.A(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload68 (.A(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload69 (.A(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload70 (.A(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload71 (.A(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload72 (.A(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload73 (.A(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload74 (.A(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload75 (.A(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload76 (.A(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload77 (.A(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload78 (.A(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload79 (.A(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload80 (.A(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload81 (.A(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload82 (.A(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload83 (.A(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload84 (.A(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload85 (.A(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload86 (.A(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload87 (.A(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload88 (.A(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload89 (.A(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload90 (.A(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload91 (.A(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload92 (.A(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload93 (.A(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload94 (.A(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload95 (.A(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload96 (.A(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload97 (.A(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload98 (.A(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload99 (.A(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkload100 (.A(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload101 (.A(clknet_leaf_27_CLK));
 sky130_fd_sc_hd__clkbuf_1 clkload102 (.A(clknet_leaf_28_CLK));
endmodule
